reg [30:0] MCODE0 [2048];
initial begin
// stateCtrl[2], addrBus[2], addrCtrl[6], regMode[5], regAXY[2], busCtrl[5], ALUCtrl[6], outBus[3]
// 00 NOP
MCODE0[0]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1]={2'b10,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[2]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[3]={2'b10,2'b00,6'b000000,5'b00011,2'b01,5'b11001,6'b100000,3'b000};// MUL207[8]: ['ALU{Y*A}', 'ALU{}->YA', 'Flags']
MCODE0[4]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b100001,3'b000};// DIV159[8-11]: ['ALU{YA/X}']
MCODE0[5]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b100001,3'b000};// ['ALU{YA/X}']
MCODE0[6]={2'b00,2'b00,6'b000000,5'b00011,2'b01,5'b11001,6'b100001,3'b000};// ['ALU{YA/X}']
MCODE0[7]={2'b10,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['ALU{}->YA', 'ALU{YA/X}', 'Flags']
// 01 TCALL 0
MCODE0[8]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']']
MCODE0[9]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[10]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[11]={2'b00,2'b10,6'b000000,5'b01101,2'b00,5'b00000,6'b000000,3'b101};// ['PCH->[SP]', 'SP--']
MCODE0[12]={2'b00,2'b10,6'b000000,5'b01101,2'b00,5'b00000,6'b000000,3'b100};// ['PCL->[SP]', 'SP--']
MCODE0[13]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[14]={2'b00,2'b11,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['[VECT]->DR']
MCODE0[15]={2'b10,2'b11,6'b000000,5'b01100,2'b00,5'b00000,6'b000000,3'b000};// ['[VECT]:DR->PC']
// 02 SET1 d.0
MCODE0[16]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[17]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[18]={2'b00,2'b01,6'b000000,5'b01011,2'b00,5'b10010,6'b010110,3'b000};// ['ALU{[AX]|01}', 'ALU{}->T']
MCODE0[19]={2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001};// ['T->[AX]']
MCODE0[20]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[21]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[22]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[23]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 03 BBS d.0
MCODE0[24]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[25]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[26]={2'b00,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['[AX]->DR']
MCODE0[27]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[28]={2'b10,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->DR', 'PC++']
MCODE0[29]={2'b00,2'b00,6'b000000,5'b01001,2'b00,5'b00000,6'b000000,3'b000};// ['PC+DR->PC']
MCODE0[30]={2'b10,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[31]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 04 OR A, d
MCODE0[32]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[33]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[34]={2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b000100,3'b000};// ['ALU{A|[AX]}', 'ALU{}->A', 'Flags']
MCODE0[35]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[36]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[37]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[38]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[39]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 05 OR A, !a
MCODE0[40]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[41]={2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'PC++']
MCODE0[42]={2'b00,2'b00,6'b001000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AH', 'PC++']
MCODE0[43]={2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b000100,3'b000};// ['ALU{A|[AX]}', 'ALU{}->A', 'Flags']
MCODE0[44]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[45]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[46]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[47]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 06 OR A, {X}
MCODE0[48]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[49]={2'b00,2'b00,6'b100101,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['X->AL', 'P->AH']
MCODE0[50]={2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b000100,3'b000};// ['ALU{A|[AX]}', 'ALU{}->A', 'Flags']
MCODE0[51]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[52]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[53]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[54]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[55]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 07 OR A, {d+X}
MCODE0[56]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[57]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[58]={2'b00,2'b00,6'b010000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['AL+X->AL']
MCODE0[59]={2'b00,2'b01,6'b110000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['[AX]->DR', 'AL+1->AL']
MCODE0[60]={2'b00,2'b01,6'b011010,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['[AX]->AH', 'DR->AL']
MCODE0[61]={2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b000100,3'b000};// ['ALU{A|[AX]}', 'ALU{}->A', 'Flags']
MCODE0[62]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[63]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 08 OR #i
MCODE0[64]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[65]={2'b10,2'b00,6'b000000,5'b00010,2'b01,5'b00000,6'b000100,3'b000};// ['ALU{A|[PC]}', 'ALU{}->A', 'Flags']
MCODE0[66]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[67]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[68]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[69]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[70]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[71]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 09 OR dd, ds
MCODE0[72]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[73]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[74]={2'b00,2'b01,6'b000000,5'b00110,2'b00,5'b00000,6'b000000,3'b000};// ['[AX]->T']
MCODE0[75]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[76]={2'b00,2'b01,6'b000000,5'b00111,2'b00,5'b01100,6'b000100,3'b000};// ['ALU{T|[AX]}', 'ALU{}->T', 'Flags']
MCODE0[77]={2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001};// ['T->[AX]']
MCODE0[78]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[79]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 0A OR1 C, m.b
MCODE0[80]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[81]={2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'PC++']
MCODE0[82]={2'b00,2'b00,6'b001000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]&1F->AH', '[PC]->DR', 'PC++']
MCODE0[83]={2'b00,2'b01,6'b000000,5'b01010,2'b00,5'b10111,6'b011001,3'b000};// ['ALU{C|[AX].b}', 'ALU{}->C']
MCODE0[84]={2'b10,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[85]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[86]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[87]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 0B ASL d
MCODE0[88]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[89]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[90]={2'b00,2'b01,6'b000000,5'b00111,2'b00,5'b00000,6'b001010,3'b000};// ['ALU{[AX]<<1}', 'ALU{}->T', 'Flags']
MCODE0[91]={2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001};// ['T->[AX]']
MCODE0[92]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[93]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[94]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[95]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 0C ASL !a
MCODE0[96]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[97]={2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'PC++']
MCODE0[98]={2'b00,2'b00,6'b001000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AH', 'PC++']
MCODE0[99]={2'b00,2'b01,6'b000000,5'b00111,2'b00,5'b00000,6'b001010,3'b000};// ['ALU{[AX]<<1}', 'ALU{}->T', 'Flags']
MCODE0[100]={2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001};// ['T->[AX]']
MCODE0[101]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[102]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[103]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 0D PUSH PSW
MCODE0[104]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[105]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[106]={2'b00,2'b10,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b011};// ['PSW->[SP]']
MCODE0[107]={2'b10,2'b10,6'b000000,5'b01101,2'b00,5'b00000,6'b000000,3'b000};// ['SP--']
MCODE0[108]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[109]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[110]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[111]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 0E TSET1 !a
MCODE0[112]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[113]={2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'PC++']
MCODE0[114]={2'b00,2'b00,6'b001000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AH', 'PC++']
MCODE0[115]={2'b00,2'b01,6'b000000,5'b00011,2'b00,5'b00000,6'b000101,3'b000};// ['ALU{[AX]}', 'Flags']
MCODE0[116]={2'b00,2'b01,6'b000000,5'b01011,2'b00,5'b00000,6'b001111,3'b000};// ['ALU{[AX]|A}', 'ALU{}->T']
MCODE0[117]={2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001};// ['T->[AX]']
MCODE0[118]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[119]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 0F BRK
MCODE0[120]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[121]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[122]={2'b00,2'b10,6'b000000,5'b01101,2'b00,5'b00000,6'b000000,3'b101};// ['PCH->[SP]', 'SP--']
MCODE0[123]={2'b00,2'b10,6'b000000,5'b01101,2'b00,5'b00000,6'b000000,3'b100};// ['PCL->[SP]', 'SP--']
MCODE0[124]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b011};// ['PSW->[SP]', 'SP--']
MCODE0[125]={2'b00,2'b00,6'b000000,5'b01111,2'b00,5'b00000,6'b000000,3'b000};// ['0->I', '1->B']
MCODE0[126]={2'b00,2'b11,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['[VECT]->DR']
MCODE0[127]={2'b10,2'b11,6'b000000,5'b01100,2'b00,5'b00000,6'b000000,3'b000};// ['[VECT]:DR->PC']
// 10 BPL
MCODE0[128]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[129]={2'b10,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->DR, 'PC++'']
MCODE0[130]={2'b00,2'b00,6'b000000,5'b01001,2'b00,5'b00000,6'b000000,3'b000};// ['PC+DR->PC']
MCODE0[131]={2'b10,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[132]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[133]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[134]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[135]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 11 TCALL 1
MCODE0[136]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[137]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[138]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[139]={2'b00,2'b10,6'b000000,5'b01101,2'b00,5'b00000,6'b000000,3'b101};// ['PCH->[SP]', 'SP--']
MCODE0[140]={2'b00,2'b10,6'b000000,5'b01101,2'b00,5'b00000,6'b000000,3'b100};// ['PCL->[SP]', 'SP--']
MCODE0[141]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[142]={2'b00,2'b11,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['[VECT]->DR']
MCODE0[143]={2'b10,2'b11,6'b000000,5'b01100,2'b00,5'b00000,6'b000000,3'b000};// ['[VECT]:DR->PC']
// 12 CLR1 d.0
MCODE0[144]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[145]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[146]={2'b00,2'b01,6'b000000,5'b01011,2'b00,5'b10010,6'b010101,3'b000};// ['ALU{[AX]&~01}', 'ALU{}->T']
MCODE0[147]={2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001};// ['T->[AX]']
MCODE0[148]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[149]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[150]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[151]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 13 BBC d.0
MCODE0[152]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[153]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[154]={2'b00,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['[AX]->DR']
MCODE0[155]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[156]={2'b10,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->DR', 'PC++']
MCODE0[157]={2'b00,2'b00,6'b000000,5'b01001,2'b00,5'b00000,6'b000000,3'b000};// ['PC+DR->PC']
MCODE0[158]={2'b10,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[159]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 14 OR A, d+X
MCODE0[160]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[161]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[162]={2'b00,2'b00,6'b010000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['AL+X->AL']
MCODE0[163]={2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b000100,3'b000};// ['ALU{A|[AX]}', 'ALU{}->A', 'Flags']
MCODE0[164]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[165]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[166]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[167]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 15 OR A, !a+X
MCODE0[168]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[169]={2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'PC++']
MCODE0[170]={2'b00,2'b00,6'b011000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AH', 'AL+X->AL', 'PC++']
MCODE0[171]={2'b00,2'b00,6'b001100,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['AH+Carry->AH']
MCODE0[172]={2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b000100,3'b000};// ['ALU{A|[AX]}', 'ALU{}->A', 'Flags']
MCODE0[173]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[174]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[175]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 16 OR A, !a+Y
MCODE0[176]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[177]={2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'PC++']
MCODE0[178]={2'b00,2'b00,6'b011001,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AH', 'AL+Y->AL', 'PC++']
MCODE0[179]={2'b00,2'b00,6'b001100,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['AH+Carry->AH']
MCODE0[180]={2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b000100,3'b000};// ['ALU{A|[AX]}', 'ALU{}->A', 'Flags']
MCODE0[181]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[182]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[183]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 17 OR A, {d}+Y
MCODE0[184]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[185]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[186]={2'b00,2'b01,6'b110000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['[AX]->DR', 'AL+1->AL']
MCODE0[187]={2'b00,2'b01,6'b011011,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['[AX]->AH', 'DR+Y->AL']
MCODE0[188]={2'b00,2'b00,6'b001100,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['AH+Carry->AH']
MCODE0[189]={2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b000100,3'b000};// ['ALU{A|[AX]}', 'ALU{}->A', 'Flags']
MCODE0[190]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[191]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 18 OR d, #i
MCODE0[192]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[193]={2'b00,2'b00,6'b000000,5'b00101,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->T', 'PC++']
MCODE0[194]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[195]={2'b00,2'b01,6'b000000,5'b00111,2'b00,5'b10000,6'b000100,3'b000};// ['ALU{T|[AX]}', 'ALU{}->T', 'Flags']
MCODE0[196]={2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001};// ['T->[AX]']
MCODE0[197]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[198]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[199]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 19 OR {X}; {Y}
MCODE0[200]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[201]={2'b00,2'b00,6'b100110,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['Y->AL', 'P->AH']
MCODE0[202]={2'b00,2'b01,6'b100101,5'b00110,2'b00,5'b00000,6'b000000,3'b000};// ['[AX]->T', 'X->AL', 'P->AH']
MCODE0[203]={2'b00,2'b01,6'b000000,5'b00111,2'b00,5'b10000,6'b000100,3'b000};// ['ALU{T|[AX]}', 'ALU{}->T', 'Flags']
MCODE0[204]={2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001};// ['T->[AX]']
MCODE0[205]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[206]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[207]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 1A DECW d
MCODE0[208]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[209]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[210]={2'b00,2'b01,6'b000000,5'b00111,2'b00,5'b10000,6'b000010,3'b000};// ['ALU{[AX]-1}', 'ALU{}->T']
MCODE0[211]={2'b00,2'b01,6'b110000,5'b00000,2'b00,5'b01100,6'b000000,3'b001};// ['T->[AX]', 'AL+1->AL']
MCODE0[212]={2'b00,2'b01,6'b000000,5'b00111,2'b00,5'b10000,6'b000001,3'b000};// ['ALU{[AX]-C}', 'ALU{}->T', 'Flags']
MCODE0[213]={2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001};// ['T->[AX]']
MCODE0[214]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[215]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 1B ASL d+X
MCODE0[216]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[217]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[218]={2'b00,2'b00,6'b010000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['AL+X->AL']
MCODE0[219]={2'b00,2'b01,6'b000000,5'b00111,2'b00,5'b00000,6'b001010,3'b000};// ['ALU{[AX]<<1}', 'ALU{}->T', 'Flags']
MCODE0[220]={2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001};// ['T->[AX]']
MCODE0[221]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[222]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[223]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 1C ASL A
MCODE0[224]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[225]={2'b10,2'b00,6'b000000,5'b00011,2'b01,5'b00001,6'b001010,3'b000};// ['ALU{A<<1}', 'ALU{}->A', 'Flags']
MCODE0[226]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[227]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[228]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[229]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[230]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[231]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 1D DEC X
MCODE0[232]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[233]={2'b10,2'b00,6'b000000,5'b00011,2'b10,5'b00101,6'b000010,3'b000};// ['ALU{X-1}', 'ALU{}->X', 'Flags']
MCODE0[234]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[235]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[236]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[237]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[238]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[239]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 1E CMP X, !a
MCODE0[240]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[241]={2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'PC++']
MCODE0[242]={2'b00,2'b00,6'b001000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AH', 'PC++']
MCODE0[243]={2'b10,2'b01,6'b000000,5'b00011,2'b00,5'b00100,6'b010011,3'b000};// ['ALU{X-[AX]}', 'Flags']
MCODE0[244]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[245]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[246]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[247]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 1F JMP [!a+X]
MCODE0[248]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[249]={2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'PC++']
MCODE0[250]={2'b00,2'b00,6'b011000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AH', 'AL+X->AL', 'PC++']
MCODE0[251]={2'b00,2'b00,6'b001100,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['AH+Carry->AH']
MCODE0[252]={2'b00,2'b01,6'b111100,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['[AX]->DR', 'AX+1->AX']
MCODE0[253]={2'b10,2'b01,6'b000000,5'b01100,2'b00,5'b00000,6'b000000,3'b000};// ['[AX]:DR->PC']
MCODE0[254]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[255]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 20 CLRP
MCODE0[256]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[257]={2'b10,2'b00,6'b000000,5'b01000,2'b00,5'b00000,6'b000000,3'b000};// ['Flags']
MCODE0[258]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[259]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[260]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[261]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[262]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[263]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 21 TCALL 2
MCODE0[264]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[265]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[266]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[267]={2'b00,2'b10,6'b000000,5'b01101,2'b00,5'b00000,6'b000000,3'b101};// ['PCH->[SP]', 'SP--']
MCODE0[268]={2'b00,2'b10,6'b000000,5'b01101,2'b00,5'b00000,6'b000000,3'b100};// ['PCL->[SP]', 'SP--']
MCODE0[269]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[270]={2'b00,2'b11,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['[VECT]->DR']
MCODE0[271]={2'b10,2'b11,6'b000000,5'b01100,2'b00,5'b00000,6'b000000,3'b000};// ['[VECT]:DR->PC']
// 22 SET1 d.1
MCODE0[272]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[273]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[274]={2'b00,2'b01,6'b000000,5'b01011,2'b00,5'b10010,6'b010110,3'b000};// ['ALU{[AX]|02}', 'ALU{}->T']
MCODE0[275]={2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001};// ['T->[AX]']
MCODE0[276]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[277]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[278]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[279]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 23 BBS d.1
MCODE0[280]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[281]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[282]={2'b00,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['[AX]->DR']
MCODE0[283]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[284]={2'b10,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->DR', 'PC++']
MCODE0[285]={2'b00,2'b00,6'b000000,5'b01001,2'b00,5'b00000,6'b000000,3'b000};// ['PC+DR->PC']
MCODE0[286]={2'b10,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[287]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 24 AND A, d
MCODE0[288]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[289]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[290]={2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b000101,3'b000};// ['ALU{[AX]}->A', 'Flags']
MCODE0[291]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[292]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[293]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[294]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[295]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 25 AND A, !a
MCODE0[296]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[297]={2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'PC++']
MCODE0[298]={2'b00,2'b00,6'b001000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AH', 'PC++']
MCODE0[299]={2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b000101,3'b000};// ['ALU{[AX]}->A', 'Flags']
MCODE0[300]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[301]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[302]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[303]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 26 AND A, {X}
MCODE0[304]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[305]={2'b00,2'b00,6'b100101,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['X->AL', 'P->AH']
MCODE0[306]={2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b000101,3'b000};// ['ALU{[AX]}->A', 'Flags']
MCODE0[307]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[308]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[309]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[310]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[311]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 27 AND A, {d+X}
MCODE0[312]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[313]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[314]={2'b00,2'b00,6'b010000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['AL+X->AL']
MCODE0[315]={2'b00,2'b01,6'b110000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['[AX]->DR', 'AL+1->AL']
MCODE0[316]={2'b00,2'b01,6'b011010,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['[AX]->AH', 'DR->AL']
MCODE0[317]={2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b000101,3'b000};// ['ALU{[AX]}->A', 'Flags']
MCODE0[318]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[319]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 28 AND #i
MCODE0[320]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[321]={2'b10,2'b00,6'b000000,5'b00010,2'b01,5'b00000,6'b000101,3'b000};// ['ALU{[PC]}->A', 'PC++', 'Flags']
MCODE0[322]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[323]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[324]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[325]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[326]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[327]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 29 AND dd, ds
MCODE0[328]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[329]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[330]={2'b00,2'b01,6'b000000,5'b00110,2'b00,5'b00000,6'b000000,3'b000};// ['[AX]->T']
MCODE0[331]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[332]={2'b00,2'b01,6'b000000,5'b00111,2'b00,5'b10000,6'b000101,3'b000};// ['ALU{[AX]}->T', 'Flags']
MCODE0[333]={2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001};// ['T->[AX]']
MCODE0[334]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[335]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 2A OR1 C, !m.b
MCODE0[336]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[337]={2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'PC++']
MCODE0[338]={2'b00,2'b00,6'b001000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]&1F->AH', 'PC++']
MCODE0[339]={2'b00,2'b01,6'b000000,5'b01010,2'b00,5'b10111,6'b011010,3'b000};// ['ALU{C|~[AX].b}', 'ALU{}->C']
MCODE0[340]={2'b10,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[341]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[342]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[343]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 2B ROL d
MCODE0[344]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[345]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[346]={2'b00,2'b01,6'b000000,5'b00111,2'b00,5'b00000,6'b001100,3'b000};// ['ALU{[AX]}->T']
MCODE0[347]={2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001};// ['T->[AX]']
MCODE0[348]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[349]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[350]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[351]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 2C ROL !a
MCODE0[352]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[353]={2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'PC++']
MCODE0[354]={2'b00,2'b00,6'b001000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AH', 'PC++']
MCODE0[355]={2'b00,2'b01,6'b000000,5'b00111,2'b00,5'b10000,6'b001100,3'b000};// ['ALU{[AX]}->T']
MCODE0[356]={2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001};// ['T->[AX]']
MCODE0[357]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[358]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[359]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 2D PUSH A
MCODE0[360]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[361]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[362]={2'b00,2'b10,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b001};// ['A->[SP]']
MCODE0[363]={2'b10,2'b10,6'b000000,5'b01101,2'b00,5'b00000,6'b000000,3'b000};// ['SP--']
MCODE0[364]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[365]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[366]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[367]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 2E CBNE d, r
MCODE0[368]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[369]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[370]={2'b00,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b010011,3'b000};// ['ALU{[AX]}']
MCODE0[371]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[372]={2'b10,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->DR', 'PC++']
MCODE0[373]={2'b00,2'b00,6'b000000,5'b01001,2'b00,5'b00000,6'b000000,3'b000};// ['PC+DR->PC']
MCODE0[374]={2'b10,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[375]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 2F BRA
MCODE0[376]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[377]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->DR', 'PC++']
MCODE0[378]={2'b00,2'b00,6'b000000,5'b01001,2'b00,5'b00000,6'b000000,3'b000};// ['PC+DR->PC']
MCODE0[379]={2'b10,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[380]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[381]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[382]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[383]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 30 BMI
MCODE0[384]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[385]={2'b10,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->DR', 'PC++']
MCODE0[386]={2'b00,2'b00,6'b000000,5'b01001,2'b00,5'b00000,6'b000000,3'b000};// ['PC+DR->PC']
MCODE0[387]={2'b10,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[388]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[389]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[390]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[391]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 31 TCALL 3
MCODE0[392]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[393]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[394]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[395]={2'b00,2'b10,6'b000000,5'b01101,2'b00,5'b00000,6'b000000,3'b101};// ['PCH->[SP]', 'SP--']
MCODE0[396]={2'b00,2'b10,6'b000000,5'b01101,2'b00,5'b00000,6'b000000,3'b100};// ['PCL->[SP]', 'SP--']
MCODE0[397]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[398]={2'b00,2'b11,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['[VECT]->DR']
MCODE0[399]={2'b10,2'b11,6'b000000,5'b01100,2'b00,5'b00000,6'b000000,3'b000};// ['[VECT]:DR->PC']
// 32 CLR1 d.1
MCODE0[400]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[401]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[402]={2'b00,2'b01,6'b000000,5'b01011,2'b00,5'b10010,6'b010101,3'b000};// ['ALU{[AX]&~02}', 'ALU{}->T']
MCODE0[403]={2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001};// ['T->[AX]']
MCODE0[404]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[405]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[406]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[407]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 33 BBC d.1
MCODE0[408]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[409]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[410]={2'b00,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['[AX]->DR']
MCODE0[411]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[412]={2'b10,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->DR', 'PC++']
MCODE0[413]={2'b00,2'b00,6'b000000,5'b01001,2'b00,5'b00000,6'b000000,3'b000};// ['PC+DR->PC']
MCODE0[414]={2'b10,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[415]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 34 AND A, d+X
MCODE0[416]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[417]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[418]={2'b00,2'b00,6'b010000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['AL+X->AL']
MCODE0[419]={2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b000101,3'b000};// ['ALU{[AX]}->A', 'Flags']
MCODE0[420]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[421]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[422]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[423]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 35 AND A, !a+X
MCODE0[424]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[425]={2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'PC++']
MCODE0[426]={2'b00,2'b00,6'b011000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AH', 'AL+X->AL', 'PC++']
MCODE0[427]={2'b00,2'b00,6'b001100,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['AH+Carry->AH']
MCODE0[428]={2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b000101,3'b000};// ['ALU{[AX]}->A', 'Flags']
MCODE0[429]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[430]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[431]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 36 AND A, !a+Y
MCODE0[432]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[433]={2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'PC++']
MCODE0[434]={2'b00,2'b00,6'b011001,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AH', 'AL+Y->AL', 'PC++']
MCODE0[435]={2'b00,2'b00,6'b001100,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['AH+Carry->AH']
MCODE0[436]={2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b000101,3'b000};// ['ALU{[AX]}->A', 'Flags']
MCODE0[437]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[438]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[439]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 37 AND A, {d}+Y
MCODE0[440]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[441]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[442]={2'b00,2'b01,6'b110000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['[AX]->DR', 'AL+1->AL']
MCODE0[443]={2'b00,2'b01,6'b011011,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['[AX]->AH', 'DR+Y->AL']
MCODE0[444]={2'b00,2'b00,6'b001100,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['AH+Carry->AH']
MCODE0[445]={2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b000101,3'b000};// ['ALU{[AX]}->A', 'Flags']
MCODE0[446]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[447]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 38 AND d, #i
MCODE0[448]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[449]={2'b00,2'b00,6'b000000,5'b00101,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->T', 'PC++']
MCODE0[450]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[451]={2'b00,2'b01,6'b000000,5'b00111,2'b00,5'b10000,6'b000101,3'b000};// ['ALU{[AX]}->T']
MCODE0[452]={2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001};// ['T->[AX]']
MCODE0[453]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[454]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[455]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 39 AND {X}; {Y}
MCODE0[456]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[457]={2'b00,2'b00,6'b100110,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['Y->AL', 'P->AH']
MCODE0[458]={2'b00,2'b01,6'b100101,5'b00110,2'b00,5'b00000,6'b000000,3'b000};// ['[AX]->T', 'X->AL', 'P->AH']
MCODE0[459]={2'b00,2'b01,6'b000000,5'b00111,2'b00,5'b10000,6'b000101,3'b000};// ['ALU{[AX]}->T']
MCODE0[460]={2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001};// ['T->[AX]']
MCODE0[461]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[462]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[463]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 3A INCW d
MCODE0[464]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[465]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[466]={2'b00,2'b01,6'b000000,5'b00111,2'b00,5'b10000,6'b000011,3'b000};// ['ALU{[AX]+1}', 'ALU{}->T']
MCODE0[467]={2'b00,2'b01,6'b110000,5'b00000,2'b00,5'b01100,6'b000000,3'b001};// ['T->[AX]', 'AL+1->AL']
MCODE0[468]={2'b00,2'b01,6'b000000,5'b00111,2'b00,5'b10000,6'b001001,3'b000};// ['ALU{[AX]+C}', 'ALU{}->T', 'Flags']
MCODE0[469]={2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001};// ['T->[AX]']
MCODE0[470]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[471]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 3B ROL d+X
MCODE0[472]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[473]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[474]={2'b00,2'b00,6'b010000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['AL+X->AL']
MCODE0[475]={2'b00,2'b01,6'b000000,5'b00111,2'b00,5'b00000,6'b001100,3'b000};// ['ALU{[AX]}->T']
MCODE0[476]={2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001};// ['T->[AX]']
MCODE0[477]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[478]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[479]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 3C ROL A
MCODE0[480]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[481]={2'b10,2'b00,6'b000000,5'b00011,2'b01,5'b00001,6'b001100,3'b000};// ['ALU{A}->A', 'Flags']
MCODE0[482]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[483]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[484]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[485]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[486]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[487]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 3D INC X
MCODE0[488]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[489]={2'b10,2'b00,6'b000000,5'b00011,2'b10,5'b00101,6'b000011,3'b000};// ['ALU{X}->X', 'Flags']
MCODE0[490]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[491]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[492]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[493]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[494]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[495]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 3E CMP X, d
MCODE0[496]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[497]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[498]={2'b10,2'b01,6'b000000,5'b00011,2'b00,5'b00100,6'b010011,3'b000};// ['ALU{X-[AX]}', 'Flags']
MCODE0[499]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[500]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[501]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[502]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[503]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 3F CALL !a
MCODE0[504]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[505]={2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'PC++']
MCODE0[506]={2'b00,2'b00,6'b001000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AH', 'PC++']
MCODE0[507]={2'b00,2'b10,6'b000000,5'b01101,2'b00,5'b00000,6'b000000,3'b101};// ['PCH->[SP]', 'SP--']
MCODE0[508]={2'b00,2'b10,6'b000000,5'b01101,2'b00,5'b00000,6'b000000,3'b100};// ['PCL->[SP]', 'SP--']
MCODE0[509]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[510]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[511]={2'b10,2'b00,6'b000000,5'b01110,2'b00,5'b00000,6'b000000,3'b000};// ['AX->PC']
// 40 SETP
MCODE0[512]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[513]={2'b10,2'b00,6'b000000,5'b01000,2'b00,5'b00000,6'b000000,3'b000};// ['Flags']
MCODE0[514]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[515]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[516]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[517]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[518]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[519]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 41 TCALL 4
MCODE0[520]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[521]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[522]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[523]={2'b00,2'b10,6'b000000,5'b01101,2'b00,5'b00000,6'b000000,3'b101};// ['PCH->[SP]', 'SP--']
MCODE0[524]={2'b00,2'b10,6'b000000,5'b01101,2'b00,5'b00000,6'b000000,3'b100};// ['PCL->[SP]', 'SP--']
MCODE0[525]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[526]={2'b00,2'b11,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['[VECT]->DR']
MCODE0[527]={2'b10,2'b11,6'b000000,5'b01100,2'b00,5'b00000,6'b000000,3'b000};// ['[VECT]:DR->PC']
// 42 SET1 d.2
MCODE0[528]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[529]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[530]={2'b00,2'b01,6'b000000,5'b01011,2'b00,5'b10010,6'b010110,3'b000};// ['ALU{[AX]|04}', 'ALU{}->T']
MCODE0[531]={2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001};// ['T->[AX]']
MCODE0[532]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[533]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[534]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[535]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 43 BBS d.2
MCODE0[536]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[537]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[538]={2'b00,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['[AX]->DR']
MCODE0[539]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[540]={2'b10,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->DR', 'PC++']
MCODE0[541]={2'b00,2'b00,6'b000000,5'b01001,2'b00,5'b00000,6'b000000,3'b000};// ['PC+DR->PC']
MCODE0[542]={2'b10,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[543]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 44 EOR A, d
MCODE0[544]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[545]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[546]={2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b000110,3'b000};// ['ALU{[AX]}->A', 'Flags']
MCODE0[547]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[548]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[549]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[550]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[551]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 45 EOR A, !a
MCODE0[552]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[553]={2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'PC++']
MCODE0[554]={2'b00,2'b00,6'b001000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AH', 'PC++']
MCODE0[555]={2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b000110,3'b000};// ['ALU{[AX]}->A', 'Flags']
MCODE0[556]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[557]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[558]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[559]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 46 EOR A, {X}
MCODE0[560]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[561]={2'b00,2'b00,6'b100101,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['X->AL', 'P->AH']
MCODE0[562]={2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b000110,3'b000};// ['ALU{[AX]}->A', 'Flags']
MCODE0[563]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[564]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[565]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[566]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[567]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 47 EOR A, {d+X}
MCODE0[568]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[569]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[570]={2'b00,2'b00,6'b010000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['AL+X->AL']
MCODE0[571]={2'b00,2'b01,6'b110000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['[AX]->DR', 'AL+1->AL']
MCODE0[572]={2'b00,2'b01,6'b011010,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['[AX]->AH', 'DR->AL']
MCODE0[573]={2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b000110,3'b000};// ['ALU{[AX]}->A', 'Flags']
MCODE0[574]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[575]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 48 EOR #i
MCODE0[576]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[577]={2'b10,2'b00,6'b000000,5'b00010,2'b01,5'b00000,6'b000110,3'b000};// ['ALU{[PC]}->A', 'PC++', 'Flags']
MCODE0[578]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[579]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[580]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[581]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[582]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[583]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 49 EOR dd, ds
MCODE0[584]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[585]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[586]={2'b00,2'b01,6'b000000,5'b00110,2'b00,5'b00000,6'b000000,3'b000};// ['[AX]->T']
MCODE0[587]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[588]={2'b00,2'b01,6'b000000,5'b00111,2'b00,5'b10000,6'b000110,3'b000};// ['ALU{[AX]}->T', 'Flags']
MCODE0[589]={2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001};// ['T->[AX]']
MCODE0[590]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[591]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 4A AND1 C, m.b
MCODE0[592]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[593]={2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'PC++']
MCODE0[594]={2'b00,2'b00,6'b001000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]&1F->AH', '[PC]->DR', 'PC++']
MCODE0[595]={2'b10,2'b01,6'b000000,5'b01010,2'b00,5'b10111,6'b010111,3'b000};// ['ALU{[AX]}->C']
MCODE0[596]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[597]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[598]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[599]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 4B LSR d
MCODE0[600]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[601]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[602]={2'b00,2'b01,6'b000000,5'b00111,2'b00,5'b00000,6'b001011,3'b000};// ['ALU{[AX]}->T']
MCODE0[603]={2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001};// ['T->[AX]']
MCODE0[604]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[605]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[606]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[607]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 4C LSR !a
MCODE0[608]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[609]={2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'PC++']
MCODE0[610]={2'b00,2'b00,6'b001000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AH', 'PC++']
MCODE0[611]={2'b00,2'b01,6'b000000,5'b00111,2'b00,5'b10000,6'b001011,3'b000};// ['ALU{[AX]}->T']
MCODE0[612]={2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001};// ['T->[AX]']
MCODE0[613]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[614]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[615]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 4D PUSH X
MCODE0[616]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[617]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[618]={2'b00,2'b10,6'b000000,5'b00000,2'b00,5'b00100,6'b000000,3'b001};// ['X->[SP]']
MCODE0[619]={2'b10,2'b10,6'b000000,5'b01101,2'b00,5'b00000,6'b000000,3'b000};// ['SP--']
MCODE0[620]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[621]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[622]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[623]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 4E TCLR1 !a
MCODE0[624]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[625]={2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'PC++']
MCODE0[626]={2'b00,2'b00,6'b001000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AH', 'PC++']
MCODE0[627]={2'b00,2'b01,6'b000000,5'b00011,2'b00,5'b00000,6'b000101,3'b000};// ['ALU{[AX]}', 'Flags']
MCODE0[628]={2'b00,2'b01,6'b000000,5'b01011,2'b00,5'b00000,6'b001110,3'b000};// ['ALU{[AX]}->T']
MCODE0[629]={2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001};// ['T->[AX]']
MCODE0[630]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[631]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 4F PCALL u
MCODE0[632]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[633]={2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'PC++']
MCODE0[634]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[635]={2'b00,2'b10,6'b000000,5'b01101,2'b00,5'b00000,6'b000000,3'b101};// ['PCH->[SP]', 'SP--']
MCODE0[636]={2'b00,2'b10,6'b000000,5'b01101,2'b00,5'b00000,6'b000000,3'b100};// ['PCL->[SP]', 'SP--']
MCODE0[637]={2'b10,2'b00,6'b000000,5'b10010,2'b00,5'b00000,6'b000000,3'b000};// ['FF:AL->PC']
MCODE0[638]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[639]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 50 BVC
MCODE0[640]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[641]={2'b10,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->DR', 'PC++']
MCODE0[642]={2'b00,2'b00,6'b000000,5'b01001,2'b00,5'b00000,6'b000000,3'b000};// ['PC+DR->PC']
MCODE0[643]={2'b10,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[644]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[645]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[646]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[647]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 51 TCALL 5
MCODE0[648]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[649]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[650]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[651]={2'b00,2'b10,6'b000000,5'b01101,2'b00,5'b00000,6'b000000,3'b101};// ['PCH->[SP]', 'SP--']
MCODE0[652]={2'b00,2'b10,6'b000000,5'b01101,2'b00,5'b00000,6'b000000,3'b100};// ['PCL->[SP]', 'SP--']
MCODE0[653]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[654]={2'b00,2'b11,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['[VECT]->DR']
MCODE0[655]={2'b10,2'b11,6'b000000,5'b01100,2'b00,5'b00000,6'b000000,3'b000};// ['[VECT]:DR->PC']
// 52 CLR1 d.2
MCODE0[656]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[657]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[658]={2'b00,2'b01,6'b000000,5'b01011,2'b00,5'b10010,6'b010101,3'b000};// ['ALU{[AX]&~04}', 'ALU{}->T']
MCODE0[659]={2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001};// ['T->[AX]']
MCODE0[660]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[661]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[662]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[663]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 53 BBC d.2
MCODE0[664]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[665]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[666]={2'b00,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['[AX]->DR']
MCODE0[667]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[668]={2'b10,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->DR', 'PC++']
MCODE0[669]={2'b00,2'b00,6'b000000,5'b01001,2'b00,5'b00000,6'b000000,3'b000};// ['PC+DR->PC']
MCODE0[670]={2'b10,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[671]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 54 EOR A, d+X
MCODE0[672]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[673]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[674]={2'b00,2'b00,6'b010000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['AL+X->AL']
MCODE0[675]={2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b000110,3'b000};// ['ALU{[AX]}->A', 'Flags']
MCODE0[676]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[677]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[678]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[679]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 55 EOR A, !a+X
MCODE0[680]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[681]={2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'PC++']
MCODE0[682]={2'b00,2'b00,6'b011000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AH', 'AL+X->AL', 'PC++']
MCODE0[683]={2'b00,2'b00,6'b001100,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['AH+Carry->AH']
MCODE0[684]={2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b000110,3'b000};// ['ALU{[AX]}->A', 'Flags']
MCODE0[685]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[686]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[687]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 56 EOR A, !a+Y
MCODE0[688]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[689]={2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'PC++']
MCODE0[690]={2'b00,2'b00,6'b011001,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AH', 'AL+X->AL', 'PC++']
MCODE0[691]={2'b00,2'b00,6'b001100,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['AH+Carry->AH']
MCODE0[692]={2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b000110,3'b000};// ['ALU{[AX]}->A', 'Flags']
MCODE0[693]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[694]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[695]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 57 EOR A, {d}+Y
MCODE0[696]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[697]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[698]={2'b00,2'b01,6'b110000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['[AX]->DR', 'AL+1->AL']
MCODE0[699]={2'b00,2'b01,6'b011011,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['[AX]->AH', 'DR+Y->AL']
MCODE0[700]={2'b00,2'b00,6'b001100,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['AH+Carry->AH']
MCODE0[701]={2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b000110,3'b000};// ['ALU{[AX]}->A', 'Flags']
MCODE0[702]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[703]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 58 EOR d, #i
MCODE0[704]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[705]={2'b00,2'b00,6'b000000,5'b00101,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->T', 'PC++']
MCODE0[706]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[707]={2'b00,2'b01,6'b000000,5'b00111,2'b00,5'b10000,6'b000110,3'b000};// ['ALU{[AX]}->T']
MCODE0[708]={2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001};// ['T->[AX]']
MCODE0[709]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[710]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[711]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 59 EOR {X}; {Y}
MCODE0[712]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[713]={2'b00,2'b00,6'b100110,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['Y->AL', 'P->AH']
MCODE0[714]={2'b00,2'b01,6'b100101,5'b00110,2'b00,5'b00000,6'b000000,3'b000};// ['[AX]->T', 'X->AL', 'P->AH']
MCODE0[715]={2'b00,2'b01,6'b000000,5'b00111,2'b00,5'b10000,6'b000110,3'b000};// ['ALU{[AX]}->T', 'Flags']
MCODE0[716]={2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001};// ['T->[AX]']
MCODE0[717]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[718]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[719]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 5A CMPW YA, d
MCODE0[720]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[721]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[722]={2'b00,2'b01,6'b000000,5'b00011,2'b00,5'b00000,6'b010011,3'b000};// ['ALU{A-[AX]}']
MCODE0[723]={2'b00,2'b01,6'b110000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['AL+1->AL']
MCODE0[724]={2'b10,2'b01,6'b000000,5'b00011,2'b00,5'b01000,6'b010000,3'b000};// ['ALU{[AX]}', 'Flags']
MCODE0[725]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[726]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[727]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 5B LSR d+X
MCODE0[728]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[729]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[730]={2'b00,2'b00,6'b010000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['AL+X->AL']
MCODE0[731]={2'b00,2'b01,6'b000000,5'b00111,2'b00,5'b00000,6'b001011,3'b000};// ['ALU{[AX]}->T']
MCODE0[732]={2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001};// ['T->[AX]']
MCODE0[733]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[734]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[735]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 5C LSR A
MCODE0[736]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[737]={2'b10,2'b00,6'b000000,5'b00011,2'b01,5'b00001,6'b001011,3'b000};// ['ALU{A}->A', 'Flags']
MCODE0[738]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[739]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[740]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[741]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[742]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[743]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 5D MOV X, A
MCODE0[744]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[745]={2'b10,2'b00,6'b000000,5'b00011,2'b10,5'b00001,6'b000000,3'b000};// ['ALU{A}->X', 'Flags']
MCODE0[746]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[747]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[748]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[749]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[750]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[751]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 5E CMP Y, !a
MCODE0[752]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[753]={2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'PC++']
MCODE0[754]={2'b00,2'b00,6'b001000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AH', 'PC++']
MCODE0[755]={2'b10,2'b01,6'b000000,5'b00011,2'b00,5'b01000,6'b010011,3'b000};// ['ALU{Y-[AX]}', 'Flags']
MCODE0[756]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[757]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[758]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[759]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 5F JMP !a
MCODE0[760]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[761]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->DR', 'PC++']
MCODE0[762]={2'b10,2'b00,6'b000000,5'b01100,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]:DR->PC']
MCODE0[763]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[764]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[765]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[766]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[767]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 60 CLRC
MCODE0[768]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[769]={2'b10,2'b00,6'b000000,5'b01000,2'b00,5'b00000,6'b000000,3'b000};// ['Flags']
MCODE0[770]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[771]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[772]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[773]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[774]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[775]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 61 TCALL 6
MCODE0[776]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[777]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[778]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[779]={2'b00,2'b10,6'b000000,5'b01101,2'b00,5'b00000,6'b000000,3'b101};// ['PCH->[SP]', 'SP--']
MCODE0[780]={2'b00,2'b10,6'b000000,5'b01101,2'b00,5'b00000,6'b000000,3'b100};// ['PCL->[SP]', 'SP--']
MCODE0[781]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[782]={2'b00,2'b11,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['[VECT]->DR']
MCODE0[783]={2'b10,2'b11,6'b000000,5'b01100,2'b00,5'b00000,6'b000000,3'b000};// ['[VECT]:DR->PC']
// 62 SET1 d.3
MCODE0[784]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[785]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[786]={2'b00,2'b01,6'b000000,5'b01011,2'b00,5'b10010,6'b010110,3'b000};// ['ALU{[AX]|08}', 'ALU{}->T']
MCODE0[787]={2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001};// ['T->[AX]']
MCODE0[788]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[789]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[790]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[791]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 63 BBS d.3
MCODE0[792]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[793]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[794]={2'b00,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['[AX]->DR']
MCODE0[795]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[796]={2'b10,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->DR', 'PC++']
MCODE0[797]={2'b00,2'b00,6'b000000,5'b01001,2'b00,5'b00000,6'b000000,3'b000};// ['PC+DR->PC']
MCODE0[798]={2'b10,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[799]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 64 CMP A, d
MCODE0[800]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[801]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[802]={2'b10,2'b01,6'b000000,5'b00011,2'b00,5'b00000,6'b010011,3'b000};// ['ALU{A-[AX]}', 'Flags']
MCODE0[803]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[804]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[805]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[806]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[807]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 65 CMP A, !a
MCODE0[808]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[809]={2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'PC++']
MCODE0[810]={2'b00,2'b00,6'b001000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AH', 'PC++']
MCODE0[811]={2'b10,2'b01,6'b000000,5'b00011,2'b00,5'b00000,6'b010011,3'b000};// ['ALU{A-[AX]}', 'Flags']
MCODE0[812]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[813]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[814]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[815]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 66 CMP A, {X}
MCODE0[816]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[817]={2'b00,2'b00,6'b100101,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['X->AL', 'P->AH']
MCODE0[818]={2'b10,2'b01,6'b000000,5'b00011,2'b00,5'b00000,6'b010011,3'b000};// ['ALU{A-[AX]}', 'Flags']
MCODE0[819]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[820]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[821]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[822]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[823]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 67 CMP A, {d+X}
MCODE0[824]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[825]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[826]={2'b00,2'b00,6'b010000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['AL+X->AL']
MCODE0[827]={2'b00,2'b01,6'b110000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['[AX]->DR', 'AL+1->AL']
MCODE0[828]={2'b00,2'b01,6'b011010,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['[AX]->AH', 'DR->AL']
MCODE0[829]={2'b10,2'b01,6'b000000,5'b00011,2'b00,5'b00000,6'b010011,3'b000};// ['ALU{A-[AX]}', 'Flags']
MCODE0[830]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[831]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 68 CMP #i
MCODE0[832]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[833]={2'b10,2'b00,6'b000000,5'b00010,2'b00,5'b00000,6'b010011,3'b000};// ['ALU{A-[PC]}', 'PC++', 'Flags']
MCODE0[834]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[835]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[836]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[837]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[838]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[839]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 69 CMP dd, ds
MCODE0[840]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[841]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[842]={2'b00,2'b01,6'b000000,5'b00110,2'b00,5'b00000,6'b000000,3'b000};// ['[AX]->T']
MCODE0[843]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[844]={2'b00,2'b01,6'b000000,5'b00111,2'b00,5'b10000,6'b010011,3'b000};// ['ALU{[AX]-T}', 'Flags']
MCODE0[845]={2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};//
MCODE0[846]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[847]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 6A AND1 C, !m.b
MCODE0[848]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[849]={2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'PC++']
MCODE0[850]={2'b00,2'b00,6'b001000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]&1F->AH', '[PC]->DR', 'PC++']
MCODE0[851]={2'b10,2'b01,6'b000000,5'b01010,2'b00,5'b10111,6'b011000,3'b000};// ['ALU{[AX]}->C']
MCODE0[852]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[853]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[854]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[855]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 6B ROR d
MCODE0[856]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[857]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[858]={2'b00,2'b01,6'b000000,5'b00111,2'b00,5'b00000,6'b001101,3'b000};// ['ALU{[AX]}->T']
MCODE0[859]={2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001};// ['T->[AX]']
MCODE0[860]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[861]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[862]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[863]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 6C ROR !a
MCODE0[864]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[865]={2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'PC++']
MCODE0[866]={2'b00,2'b00,6'b001000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AH', 'PC++']
MCODE0[867]={2'b00,2'b01,6'b000000,5'b00111,2'b00,5'b10000,6'b001101,3'b000};// ['ALU{[AX]}->T']
MCODE0[868]={2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001};// ['T->[AX]']
MCODE0[869]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[870]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[871]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 6D PUSH Y
MCODE0[872]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[873]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[874]={2'b00,2'b10,6'b000000,5'b00000,2'b00,5'b01000,6'b000000,3'b001};// ['Y->[SP]']
MCODE0[875]={2'b10,2'b10,6'b000000,5'b01101,2'b00,5'b00000,6'b000000,3'b000};// ['SP--']
MCODE0[876]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[877]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[878]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[879]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 6E DBNZ d, r
MCODE0[880]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[881]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[882]={2'b00,2'b01,6'b000000,5'b00111,2'b00,5'b10000,6'b000010,3'b000};// ['ALU{[AX]}->T']
MCODE0[883]={2'b00,2'b01,6'b000000,5'b00000,2'b00,5'b01101,6'b000000,3'b001};// ['T->[AX]']
MCODE0[884]={2'b10,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->DR', 'PC++']
MCODE0[885]={2'b00,2'b00,6'b000000,5'b01001,2'b00,5'b00000,6'b000000,3'b000};// ['PC+DR->PC']
MCODE0[886]={2'b10,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[887]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 6F RET
MCODE0[888]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[889]={2'b00,2'b00,6'b000000,5'b10000,2'b00,5'b00000,6'b000000,3'b000};// ['SP++']
MCODE0[890]={2'b00,2'b10,6'b000000,5'b10000,2'b00,5'b00000,6'b000000,3'b000};// ['[SP]->DR', 'SP++']
MCODE0[891]={2'b00,2'b10,6'b000000,5'b01100,2'b00,5'b00000,6'b000000,3'b000};// ['[SP]:DR->PC']
MCODE0[892]={2'b10,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[893]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[894]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[895]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 70 BVS
MCODE0[896]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[897]={2'b10,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->DR', 'PC++']
MCODE0[898]={2'b00,2'b00,6'b000000,5'b01001,2'b00,5'b00000,6'b000000,3'b000};// ['PC+DR->PC']
MCODE0[899]={2'b10,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[900]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[901]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[902]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[903]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 71 TCALL 7
MCODE0[904]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[905]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[906]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[907]={2'b00,2'b10,6'b000000,5'b01101,2'b00,5'b00000,6'b000000,3'b101};// ['PCH->[SP]', 'SP--']
MCODE0[908]={2'b00,2'b10,6'b000000,5'b01101,2'b00,5'b00000,6'b000000,3'b100};// ['PCL->[SP]', 'SP--']
MCODE0[909]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[910]={2'b00,2'b11,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['[VECT]->DR']
MCODE0[911]={2'b10,2'b11,6'b000000,5'b01100,2'b00,5'b00000,6'b000000,3'b000};// ['[VECT]:DR->PC']
// 72 CLR1 d.3
MCODE0[912]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[913]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[914]={2'b00,2'b01,6'b000000,5'b01011,2'b00,5'b10010,6'b010101,3'b000};// ['ALU{[AX]&~08}', 'ALU{}->T']
MCODE0[915]={2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001};// ['T->[AX]']
MCODE0[916]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[917]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[918]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[919]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 73 BBC d.3
MCODE0[920]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[921]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[922]={2'b00,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['[AX]->DR']
MCODE0[923]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[924]={2'b10,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->DR', 'PC++']
MCODE0[925]={2'b00,2'b00,6'b000000,5'b01001,2'b00,5'b00000,6'b000000,3'b000};// ['PC+DR->PC']
MCODE0[926]={2'b10,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[927]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 74 CMP A, d+X
MCODE0[928]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[929]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[930]={2'b00,2'b00,6'b010000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['AL+X->AL']
MCODE0[931]={2'b10,2'b01,6'b000000,5'b00011,2'b00,5'b00000,6'b010011,3'b000};// ['ALU{A-[AX]}', 'Flags']
MCODE0[932]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[933]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[934]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[935]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 75 CMP A, !a+X
MCODE0[936]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[937]={2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'PC++']
MCODE0[938]={2'b00,2'b00,6'b011000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AH', 'AL+X->AL', 'PC++']
MCODE0[939]={2'b00,2'b00,6'b001100,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['AH+Carry->AH']
MCODE0[940]={2'b10,2'b01,6'b000000,5'b00011,2'b00,5'b00000,6'b010011,3'b000};// ['ALU{A-[AX]}', 'Flags']
MCODE0[941]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[942]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[943]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 76 CMP A, !a+Y
MCODE0[944]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[945]={2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'PC++']
MCODE0[946]={2'b00,2'b00,6'b011001,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AH', 'AL+X->AL', 'PC++']
MCODE0[947]={2'b00,2'b00,6'b001100,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['AH+Carry->AH']
MCODE0[948]={2'b10,2'b01,6'b000000,5'b00011,2'b00,5'b00000,6'b010011,3'b000};// ['ALU{A-[AX]}', 'Flags']
MCODE0[949]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[950]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[951]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 77 CMP A, {d}+Y
MCODE0[952]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[953]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[954]={2'b00,2'b01,6'b110000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['[AX]->DR', 'AL+1->AL']
MCODE0[955]={2'b00,2'b01,6'b011011,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['[AX]->AH', 'DR+Y->AL']
MCODE0[956]={2'b00,2'b00,6'b001100,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['AH+Carry->AH']
MCODE0[957]={2'b10,2'b01,6'b000000,5'b00011,2'b00,5'b00000,6'b010011,3'b000};// ['ALU{A-[AX]}', 'Flags']
MCODE0[958]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[959]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 78 CMP d, #i
MCODE0[960]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[961]={2'b00,2'b00,6'b000000,5'b00101,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->T', 'PC++']
MCODE0[962]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[963]={2'b00,2'b01,6'b000000,5'b00111,2'b00,5'b10000,6'b010011,3'b000};// ['ALU{[AX]-T}', 'Flags']
MCODE0[964]={2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};//
MCODE0[965]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[966]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[967]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 79 CMP {X}; {Y}
MCODE0[968]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[969]={2'b00,2'b00,6'b100110,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['Y->AL', 'P->AH']
MCODE0[970]={2'b00,2'b01,6'b100101,5'b00110,2'b00,5'b00000,6'b000000,3'b000};// ['[AX]->T', 'X->AL', 'P->AH']
MCODE0[971]={2'b00,2'b01,6'b000000,5'b00111,2'b00,5'b10000,6'b010011,3'b000};// ['ALU{[AX]-T}', 'Flags']
MCODE0[972]={2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};//
MCODE0[973]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[974]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[975]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 7A ADDW YA, d
MCODE0[976]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[977]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[978]={2'b00,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b010001,3'b000};// ['ALU{[AX]}->A']
MCODE0[979]={2'b00,2'b00,6'b110000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['AL+1->AL']
MCODE0[980]={2'b10,2'b01,6'b000000,5'b00011,2'b11,5'b01000,6'b010010,3'b000};// ['ALU{[AX]}->Y']
MCODE0[981]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[982]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[983]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 7B ROR d+X
MCODE0[984]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[985]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[986]={2'b00,2'b00,6'b010000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['AL+X->AL']
MCODE0[987]={2'b00,2'b01,6'b000000,5'b00111,2'b00,5'b00000,6'b001101,3'b000};// ['ALU{[AX]}->T']
MCODE0[988]={2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001};// ['T->[AX]']
MCODE0[989]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[990]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[991]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 7C ROR A
MCODE0[992]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[993]={2'b10,2'b00,6'b000000,5'b00011,2'b01,5'b00001,6'b001101,3'b000};// ['ALU{A}->A', 'Flags']
MCODE0[994]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[995]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[996]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[997]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[998]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[999]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 7D MOV A, X
MCODE0[1000]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1001]={2'b10,2'b00,6'b000000,5'b00011,2'b01,5'b00101,6'b000000,3'b000};// ['ALU{X}->A', 'Flags']
MCODE0[1002]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1003]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1004]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1005]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1006]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1007]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 7E CMP Y, d
MCODE0[1008]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1009]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[1010]={2'b10,2'b01,6'b000000,5'b00011,2'b00,5'b01000,6'b010011,3'b000};// ['ALU{Y-[AX]}', 'Flags']
MCODE0[1011]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1012]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1013]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1014]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1015]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 7F RETI
MCODE0[1016]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1017]={2'b00,2'b00,6'b000000,5'b10000,2'b00,5'b00000,6'b000000,3'b000};// ['SP++']
MCODE0[1018]={2'b00,2'b10,6'b000000,5'b10001,2'b00,5'b00000,6'b000000,3'b000};// ['[SP]->PSW']
MCODE0[1019]={2'b00,2'b00,6'b000000,5'b10000,2'b00,5'b00000,6'b000000,3'b000};// ['SP++']
MCODE0[1020]={2'b00,2'b10,6'b000000,5'b10000,2'b00,5'b00000,6'b000000,3'b000};// ['[SP]->DR', 'SP++']
MCODE0[1021]={2'b10,2'b10,6'b000000,5'b01100,2'b00,5'b00000,6'b000000,3'b000};// ['[SP]:DR->PC']
MCODE0[1022]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1023]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 80 SETC
MCODE0[1024]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1025]={2'b10,2'b00,6'b000000,5'b01000,2'b00,5'b00000,6'b000000,3'b000};// ['Flags']
MCODE0[1026]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1027]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1028]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1029]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1030]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1031]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 81 TCALL 8
MCODE0[1032]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1033]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[1034]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[1035]={2'b00,2'b10,6'b000000,5'b01101,2'b00,5'b00000,6'b000000,3'b101};// ['PCH->[SP]', 'SP--']
MCODE0[1036]={2'b00,2'b10,6'b000000,5'b01101,2'b00,5'b00000,6'b000000,3'b100};// ['PCL->[SP]', 'SP--']
MCODE0[1037]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[1038]={2'b00,2'b11,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['[VECT]->DR']
MCODE0[1039]={2'b10,2'b11,6'b000000,5'b01100,2'b00,5'b00000,6'b000000,3'b000};// ['[VECT]:DR->PC']
// 82 SET1 d.4
MCODE0[1040]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1041]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[1042]={2'b00,2'b01,6'b000000,5'b01011,2'b00,5'b10010,6'b010110,3'b000};// ['ALU{[AX]|10}', 'ALU{}->T']
MCODE0[1043]={2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001};// ['T->[AX]']
MCODE0[1044]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1045]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1046]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1047]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 83 BBS d.4
MCODE0[1048]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1049]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[1050]={2'b00,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['[AX]->DR']
MCODE0[1051]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[1052]={2'b10,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->DR', 'PC++']
MCODE0[1053]={2'b00,2'b00,6'b000000,5'b01001,2'b00,5'b00000,6'b000000,3'b000};// ['PC+DR->PC']
MCODE0[1054]={2'b10,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[1055]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 84 ADC A, d
MCODE0[1056]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1057]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[1058]={2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b000111,3'b000};// ['ALU{[AX]}->A', 'Flags']
MCODE0[1059]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1060]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1061]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1062]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1063]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 85 ADC A, !a
MCODE0[1064]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1065]={2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'PC++']
MCODE0[1066]={2'b00,2'b00,6'b001000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AH', 'PC++']
MCODE0[1067]={2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b000111,3'b000};// ['ALU{[AX]}->A', 'Flags']
MCODE0[1068]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1069]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1070]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1071]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 86 ADC A, {X}
MCODE0[1072]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1073]={2'b00,2'b00,6'b100101,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['X->AL', 'P->AH']
MCODE0[1074]={2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b000111,3'b000};// ['ALU{[AX]}->A', 'Flags']
MCODE0[1075]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1076]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1077]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1078]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1079]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 87 ADC A, {d+X}
MCODE0[1080]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1081]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[1082]={2'b00,2'b00,6'b010000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['AL+X->AL']
MCODE0[1083]={2'b00,2'b01,6'b110000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['[AX]->DR', 'AL+1->AL']
MCODE0[1084]={2'b00,2'b01,6'b011010,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['[AX]->AH', 'DR->AL']
MCODE0[1085]={2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b000111,3'b000};// ['ALU{[AX]}->A', 'Flags']
MCODE0[1086]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1087]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 88 ADC #i
MCODE0[1088]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1089]={2'b10,2'b00,6'b000000,5'b00010,2'b01,5'b00000,6'b000111,3'b000};// ['ALU{[PC]}->A', 'PC++', 'Flags']
MCODE0[1090]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1091]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1092]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1093]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1094]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1095]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 89 ADC dd, ds
MCODE0[1096]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1097]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[1098]={2'b00,2'b01,6'b000000,5'b00110,2'b00,5'b00000,6'b000000,3'b000};// ['[AX]->T']
MCODE0[1099]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[1100]={2'b00,2'b01,6'b000000,5'b00111,2'b00,5'b10000,6'b000111,3'b000};// ['ALU{[AX]}->T', 'Flags']
MCODE0[1101]={2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001};// ['T->[AX]']
MCODE0[1102]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1103]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 8A EOR1 C, m.b
MCODE0[1104]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1105]={2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'PC++']
MCODE0[1106]={2'b00,2'b00,6'b001000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]&1F->AH', '[PC]->DR', 'PC++']
MCODE0[1107]={2'b10,2'b01,6'b000000,5'b01010,2'b00,5'b10111,6'b011011,3'b000};// ['ALU{[AX]}->C']
MCODE0[1108]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1109]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1110]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1111]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 8B DEC d
MCODE0[1112]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1113]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[1114]={2'b00,2'b01,6'b000000,5'b00111,2'b00,5'b10000,6'b000010,3'b000};// ['ALU{[AX]-1}', 'ALU{}->T', 'Flags']
MCODE0[1115]={2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001};// ['T->[AX]']
MCODE0[1116]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1117]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1118]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1119]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 8C DEC !a
MCODE0[1120]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1121]={2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'PC++']
MCODE0[1122]={2'b00,2'b00,6'b001000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AH', 'PC++']
MCODE0[1123]={2'b00,2'b01,6'b000000,5'b00111,2'b00,5'b10000,6'b000010,3'b000};// ['ALU{[AX]-1}', 'ALU{}->T', 'Flags']
MCODE0[1124]={2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001};// ['T->[AX]']
MCODE0[1125]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1126]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1127]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 8D MOV Y, #i
MCODE0[1128]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1129]={2'b10,2'b00,6'b000000,5'b00010,2'b11,5'b00000,6'b000000,3'b000};// ['ALU{[PC]}->Y', 'PC++', 'Flags']
MCODE0[1130]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1131]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1132]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1133]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1134]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1135]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 8E POP PSW
MCODE0[1136]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1137]={2'b00,2'b00,6'b000000,5'b10000,2'b00,5'b00000,6'b000000,3'b000};// ['SP++']
MCODE0[1138]={2'b10,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[1139]={2'b00,2'b10,6'b000000,5'b10001,2'b00,5'b00000,6'b000000,3'b000};// ['[SP]->PSW']
MCODE0[1140]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1141]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1142]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1143]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 8F MOV d, #i
MCODE0[1144]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1145]={2'b00,2'b00,6'b000000,5'b00101,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->T', 'PC++']
MCODE0[1146]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[1147]={2'b00,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['[AX]']
MCODE0[1148]={2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001};// ['T->[AX]']
MCODE0[1149]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1150]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1151]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 90 BCC
MCODE0[1152]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1153]={2'b10,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->DR', 'PC++']
MCODE0[1154]={2'b00,2'b00,6'b000000,5'b01001,2'b00,5'b00000,6'b000000,3'b000};// ['PC+DR->PC']
MCODE0[1155]={2'b10,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[1156]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1157]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1158]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1159]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 91 TCALL 9
MCODE0[1160]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1161]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[1162]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[1163]={2'b00,2'b10,6'b000000,5'b01101,2'b00,5'b00000,6'b000000,3'b101};// ['PCH->[SP]', 'SP--']
MCODE0[1164]={2'b00,2'b10,6'b000000,5'b01101,2'b00,5'b00000,6'b000000,3'b100};// ['PCL->[SP]', 'SP--']
MCODE0[1165]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[1166]={2'b00,2'b11,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['[VECT]->DR']
MCODE0[1167]={2'b10,2'b11,6'b000000,5'b01100,2'b00,5'b00000,6'b000000,3'b000};// ['[VECT]:DR->PC']
// 92 CLR1 d.4
MCODE0[1168]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1169]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[1170]={2'b00,2'b01,6'b000000,5'b01011,2'b00,5'b10010,6'b010101,3'b000};// ['ALU{[AX]&~10}', 'ALU{}->T']
MCODE0[1171]={2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001};// ['T->[AX]']
MCODE0[1172]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1173]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1174]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1175]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 93 BBC d.4
MCODE0[1176]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1177]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[1178]={2'b00,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['[AX]->DR']
MCODE0[1179]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[1180]={2'b10,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->DR', 'PC++']
MCODE0[1181]={2'b00,2'b00,6'b000000,5'b01001,2'b00,5'b00000,6'b000000,3'b000};// ['PC+DR->PC']
MCODE0[1182]={2'b10,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[1183]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 94 ADC A, d+X
MCODE0[1184]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1185]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[1186]={2'b00,2'b00,6'b010000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['AL+X->AL']
MCODE0[1187]={2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b000111,3'b000};// ['ALU{[AX]}->A', 'Flags']
MCODE0[1188]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1189]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1190]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1191]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 95 ADC A, !a+X
MCODE0[1192]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1193]={2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'PC++']
MCODE0[1194]={2'b00,2'b00,6'b011000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AH', 'AL+X->AL', 'PC++']
MCODE0[1195]={2'b00,2'b00,6'b001100,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['AH+Carry->AH']
MCODE0[1196]={2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b000111,3'b000};// ['ALU{[AX]}->A', 'Flags']
MCODE0[1197]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1198]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1199]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 96 ADC A, !a+Y
MCODE0[1200]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1201]={2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'PC++']
MCODE0[1202]={2'b00,2'b00,6'b011001,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AH', 'AL+X->AL', 'PC++']
MCODE0[1203]={2'b00,2'b00,6'b001100,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['AH+Carry->AH']
MCODE0[1204]={2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b000111,3'b000};// ['ALU{[AX]}->A', 'Flags']
MCODE0[1205]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1206]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1207]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 97 ADC A, {d}+Y
MCODE0[1208]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1209]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[1210]={2'b00,2'b01,6'b110000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['[AX]->DR', 'AL+1->AL']
MCODE0[1211]={2'b00,2'b01,6'b011011,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['[AX]->AH', 'DR+Y->AL']
MCODE0[1212]={2'b00,2'b00,6'b001100,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['AH+Carry->AH']
MCODE0[1213]={2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b000111,3'b000};// ['ALU{[AX]}->A', 'Flags']
MCODE0[1214]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1215]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 98 ADC d, #i
MCODE0[1216]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1217]={2'b00,2'b00,6'b000000,5'b00101,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->T', 'PC++']
MCODE0[1218]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[1219]={2'b00,2'b01,6'b000000,5'b00111,2'b00,5'b10000,6'b000111,3'b000};// ['ALU{[AX]}->T']
MCODE0[1220]={2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001};// ['T->[AX]']
MCODE0[1221]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1222]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1223]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 99 ADC {X}; {Y}
MCODE0[1224]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1225]={2'b00,2'b00,6'b100110,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['Y->AL', 'P->AH']
MCODE0[1226]={2'b00,2'b01,6'b100101,5'b00110,2'b00,5'b00000,6'b000000,3'b000};// ['[AX]->T', 'X->AL', 'P->AH']
MCODE0[1227]={2'b00,2'b01,6'b000000,5'b00111,2'b00,5'b10000,6'b000111,3'b000};// ['ALU{[AX]}->T']
MCODE0[1228]={2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001};// ['T->[AX]']
MCODE0[1229]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1230]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1231]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 9A SUBW YA, d
MCODE0[1232]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1233]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[1234]={2'b00,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b010011,3'b000};// ['ALU{[AX]}->A']
MCODE0[1235]={2'b00,2'b01,6'b110000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['AL+1->AL']
MCODE0[1236]={2'b10,2'b01,6'b000000,5'b00011,2'b11,5'b01000,6'b010100,3'b000};// ['ALU{[AX]}->Y']
MCODE0[1237]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1238]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1239]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 9B DEC d+X
MCODE0[1240]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1241]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[1242]={2'b00,2'b00,6'b010000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['AL+X->AL']
MCODE0[1243]={2'b00,2'b01,6'b000000,5'b00111,2'b00,5'b10000,6'b000010,3'b000};// ['ALU{[AX]-1}', 'ALU{}->T', 'Flags']
MCODE0[1244]={2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001};// ['T->[AX]']
MCODE0[1245]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1246]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1247]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 9C DEC A
MCODE0[1248]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1249]={2'b10,2'b00,6'b000000,5'b00011,2'b01,5'b00001,6'b000010,3'b000};// ['ALU{A-1}', 'ALU{}->A', 'Flags']
MCODE0[1250]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1251]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1252]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1253]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1254]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1255]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 9D MOV X, SP
MCODE0[1256]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1257]={2'b10,2'b00,6'b000000,5'b00011,2'b10,5'b11101,6'b000000,3'b000};// ['ALU{SP}->X', 'Flags']
MCODE0[1258]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1259]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1260]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1261]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1262]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1263]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// 9E DIV YA, X
MCODE0[1264]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1265]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b100001,3'b000};// ['ALU{YA/X}']
MCODE0[1266]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b100001,3'b000};// ['ALU{YA/X}']
MCODE0[1267]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b100001,3'b000};// ['ALU{YA/X}']
MCODE0[1268]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b100001,3'b000};// ['ALU{YA/X}']
MCODE0[1269]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b100001,3'b000};// ['ALU{YA/X}']
MCODE0[1270]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b100001,3'b000};// ['ALU{YA/X}']
MCODE0[1271]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b100001,3'b000};// ['ALU{YA/X}']
// 9F XCN
MCODE0[1272]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1273]={2'b00,2'b00,6'b000000,5'b00011,2'b01,5'b00001,6'b011101,3'b000};// ['ALU{A}->A', 'Flags']
MCODE0[1274]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};
MCODE0[1275]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};
MCODE0[1276]={2'b10,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};
MCODE0[1277]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1278]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1279]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
//A0 EI
MCODE0[1280]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1281]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[1282]={2'b10,2'b00,6'b000000,5'b01000,2'b00,5'b00000,6'b000000,3'b000};// ['Flags']
MCODE0[1283]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1284]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1285]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1286]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1287]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// A1 TCALL 10
MCODE0[1288]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1289]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[1290]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[1291]={2'b00,2'b10,6'b000000,5'b01101,2'b00,5'b00000,6'b000000,3'b101};// ['PCH->[SP]', 'SP--']
MCODE0[1292]={2'b00,2'b10,6'b000000,5'b01101,2'b00,5'b00000,6'b000000,3'b100};// ['PCL->[SP]', 'SP--']
MCODE0[1293]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[1294]={2'b00,2'b11,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['[VECT]->DR']
MCODE0[1295]={2'b10,2'b11,6'b000000,5'b01100,2'b00,5'b00000,6'b000000,3'b000};// ['[VECT]:DR->PC']
// A2 SET1 d.5
MCODE0[1296]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1297]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[1298]={2'b00,2'b01,6'b000000,5'b01011,2'b00,5'b10010,6'b010110,3'b000};// ['ALU{[AX]|20}', 'ALU{}->T']
MCODE0[1299]={2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001};// ['T->[AX]']
MCODE0[1300]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1301]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1302]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1303]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// A3 BBS d.5
MCODE0[1304]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1305]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[1306]={2'b00,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['[AX]->DR']
MCODE0[1307]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[1308]={2'b10,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->DR', 'PC++']
MCODE0[1309]={2'b00,2'b00,6'b000000,5'b01001,2'b00,5'b00000,6'b000000,3'b000};// ['PC+DR->PC']
MCODE0[1310]={2'b10,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[1311]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// A4 SBC A, d
MCODE0[1312]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1313]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[1314]={2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b001000,3'b000};// ['ALU{[AX]}->A', 'Flags']
MCODE0[1315]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1316]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1317]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1318]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1319]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// A5 SBC A, !a
MCODE0[1320]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1321]={2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'PC++']
MCODE0[1322]={2'b00,2'b00,6'b001000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AH', 'PC++']
MCODE0[1323]={2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b001000,3'b000};// ['ALU{[AX]}->A', 'Flags']
MCODE0[1324]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1325]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1326]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1327]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// A6 SBC A, {X}
MCODE0[1328]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1329]={2'b00,2'b00,6'b100101,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['X->AL', 'P->AH']
MCODE0[1330]={2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b001000,3'b000};// ['ALU{[AX]}->A', 'Flags']
MCODE0[1331]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1332]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1333]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1334]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1335]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// A7 SBC A, {d+X}
MCODE0[1336]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1337]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[1338]={2'b00,2'b00,6'b010000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['AL+X->AL']
MCODE0[1339]={2'b00,2'b01,6'b110000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['[AX]->DR', 'AL+1->AL']
MCODE0[1340]={2'b00,2'b01,6'b011010,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['[AX]->AH', 'DR->AL']
MCODE0[1341]={2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b001000,3'b000};// ['ALU{[AX]}->A', 'Flags']
MCODE0[1342]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1343]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// A8 SBC #i
MCODE0[1344]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1345]={2'b10,2'b00,6'b000000,5'b00010,2'b01,5'b00000,6'b001000,3'b000};// ['ALU{[PC]}->A', 'PC++', 'Flags']
MCODE0[1346]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1347]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1348]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1349]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1350]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1351]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// A9 SBC dd, ds
MCODE0[1352]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1353]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[1354]={2'b00,2'b01,6'b000000,5'b00110,2'b00,5'b00000,6'b000000,3'b000};// ['[AX]->T']
MCODE0[1355]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[1356]={2'b00,2'b01,6'b000000,5'b00111,2'b00,5'b10000,6'b001000,3'b000};// ['ALU{[AX]}->T', 'Flags']
MCODE0[1357]={2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001};// ['T->[AX]']
MCODE0[1358]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1359]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// AA MOV1 C, m.b
MCODE0[1360]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1361]={2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'PC++']
MCODE0[1362]={2'b00,2'b00,6'b001000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]&1F->AH', '[PC]->DR', 'PC++']
MCODE0[1363]={2'b10,2'b01,6'b000000,5'b01010,2'b00,5'b00011,6'b000000,3'b000};// ['ALU{[AX]}->C']
MCODE0[1364]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1365]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1366]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1367]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// AB INC d
MCODE0[1368]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1369]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[1370]={2'b00,2'b01,6'b000000,5'b00111,2'b00,5'b10000,6'b000011,3'b000};// ['ALU{[AX]}->T']
MCODE0[1371]={2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001};// ['T->[AX]']
MCODE0[1372]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1373]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1374]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1375]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// AC INC !a
MCODE0[1376]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1377]={2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'PC++']
MCODE0[1378]={2'b00,2'b00,6'b001000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AH', 'PC++']
MCODE0[1379]={2'b00,2'b01,6'b000000,5'b00111,2'b00,5'b10000,6'b000011,3'b000};// ['ALU{[AX]}->T']
MCODE0[1380]={2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001};// ['T->[AX]']
MCODE0[1381]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1382]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1383]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// AD CMP Y, #i
MCODE0[1384]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1385]={2'b10,2'b00,6'b000000,5'b00010,2'b00,5'b01000,6'b010011,3'b000};// ['ALU{Y-[PC]}; 'PC++', 'Flags']
MCODE0[1386]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1387]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1388]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1389]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1390]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1391]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// AE POP A
MCODE0[1392]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1393]={2'b00,2'b00,6'b000000,5'b10000,2'b00,5'b00000,6'b000000,3'b000};// ['SP++']
MCODE0[1394]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[1395]={2'b10,2'b10,6'b000000,5'b00000,2'b01,5'b00000,6'b000000,3'b000};// ['[SP]->A']
MCODE0[1396]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1397]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1398]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1399]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// AF MOV {X}+, A
MCODE0[1400]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1401]={2'b00,2'b00,6'b100101,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['X->AL', 'P->AH']
MCODE0[1402]={2'b00,2'b00,6'b000000,5'b00000,2'b10,5'b00101,6'b000011,3'b000};// ['X++']
MCODE0[1403]={2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b001};// ['A->[AX]']
MCODE0[1404]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1405]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1406]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1407]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// B0 BCS
MCODE0[1408]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1409]={2'b10,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->DR', 'PC++']
MCODE0[1410]={2'b00,2'b00,6'b000000,5'b01001,2'b00,5'b00000,6'b000000,3'b000};// ['PC+DR->PC']
MCODE0[1411]={2'b10,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[1412]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1413]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1414]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1415]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// B1 TCALL 11
MCODE0[1416]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1417]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[1418]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[1419]={2'b00,2'b10,6'b000000,5'b01101,2'b00,5'b00000,6'b000000,3'b101};// ['PCH->[SP]', 'SP--']
MCODE0[1420]={2'b00,2'b10,6'b000000,5'b01101,2'b00,5'b00000,6'b000000,3'b100};// ['PCL->[SP]', 'SP--']
MCODE0[1421]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[1422]={2'b00,2'b11,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['[VECT]->DR']
MCODE0[1423]={2'b10,2'b11,6'b000000,5'b01100,2'b00,5'b00000,6'b000000,3'b000};// ['[VECT]:DR->PC']
// B2 CLR1 d.5
MCODE0[1424]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1425]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[1426]={2'b00,2'b01,6'b000000,5'b01011,2'b00,5'b10010,6'b010101,3'b000};// ['ALU{[AX]&~20}', 'ALU{}->T']
MCODE0[1427]={2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001};// ['T->[AX]']
MCODE0[1428]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1429]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1430]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1431]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// B3 BBC d.5
MCODE0[1432]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1433]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[1434]={2'b00,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['[AX]->DR']
MCODE0[1435]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[1436]={2'b10,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->DR', 'PC++']
MCODE0[1437]={2'b00,2'b00,6'b000000,5'b01001,2'b00,5'b00000,6'b000000,3'b000};// ['PC+DR->PC']
MCODE0[1438]={2'b10,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[1439]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// B4 SBC A, d+X
MCODE0[1440]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1441]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[1442]={2'b00,2'b00,6'b010000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['AL+X->AL']
MCODE0[1443]={2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b001000,3'b000};// ['ALU{[AX]}->A', 'Flags']
MCODE0[1444]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1445]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1446]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1447]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// B5 SBC A, !a+X
MCODE0[1448]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1449]={2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'PC++']
MCODE0[1450]={2'b00,2'b00,6'b011000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AH', 'AL+X->AL', 'PC++']
MCODE0[1451]={2'b00,2'b00,6'b001100,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['AH+Carry->AH']
MCODE0[1452]={2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b001000,3'b000};// ['ALU{[AX]}->A', 'Flags']
MCODE0[1453]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1454]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1455]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// B6 SBC A, !a+Y
MCODE0[1456]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1457]={2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'PC++']
MCODE0[1458]={2'b00,2'b00,6'b011001,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AH', 'AL+X->AL', 'PC++']
MCODE0[1459]={2'b00,2'b00,6'b001100,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['AH+Carry->AH']
MCODE0[1460]={2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b001000,3'b000};// ['ALU{[AX]}->A', 'Flags']
MCODE0[1461]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1462]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1463]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// B7 SBC A, {d}+Y
MCODE0[1464]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1465]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[1466]={2'b00,2'b01,6'b110000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['[AX]->DR', 'AL+1->AL']
MCODE0[1467]={2'b00,2'b01,6'b011011,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['[AX]->AH', 'DR+Y->AL']
MCODE0[1468]={2'b00,2'b00,6'b001100,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['AH+Carry->AH']
MCODE0[1469]={2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b001000,3'b000};// ['ALU{[AX]}->A', 'Flags']
MCODE0[1470]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1471]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// B8 SBC d, #i
MCODE0[1472]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1473]={2'b00,2'b00,6'b000000,5'b00101,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->T', 'PC++']
MCODE0[1474]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[1475]={2'b00,2'b01,6'b000000,5'b00111,2'b00,5'b10000,6'b001000,3'b000};// ['ALU{[AX]}->T']
MCODE0[1476]={2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001};// ['T->[AX]']
MCODE0[1477]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1478]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1479]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// B9 SBC {X}; {Y}
MCODE0[1480]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1481]={2'b00,2'b00,6'b100110,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['Y->AL', 'P->AH']
MCODE0[1482]={2'b00,2'b01,6'b100101,5'b00110,2'b00,5'b00000,6'b000000,3'b000};// ['[AX]->T', 'X->AL', 'P->AH']
MCODE0[1483]={2'b00,2'b01,6'b000000,5'b00111,2'b00,5'b10000,6'b001000,3'b000};// ['ALU{[AX]}->T']
MCODE0[1484]={2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001};// ['T->[AX]']
MCODE0[1485]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1486]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1487]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// BA MOV YA, d
MCODE0[1488]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1489]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[1490]={2'b00,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b000000,3'b000};// ['ALU{[AX]}->A', 'Flags']
MCODE0[1491]={2'b00,2'b00,6'b110000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['AL+1->AL']
MCODE0[1492]={2'b10,2'b01,6'b000000,5'b00011,2'b11,5'b00000,6'b000000,3'b000};// ['ALU{[AX]}->Y', 'Flags']
MCODE0[1493]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1494]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1495]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// BB INC d+X
MCODE0[1496]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1497]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[1498]={2'b00,2'b00,6'b010000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['AL+X->AL']
MCODE0[1499]={2'b00,2'b01,6'b000000,5'b00111,2'b00,5'b10000,6'b000011,3'b000};// ['ALU{[AX]}->T']
MCODE0[1500]={2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001};// ['T->[AX]']
MCODE0[1501]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1502]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1503]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// BC INC A
MCODE0[1504]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1505]={2'b10,2'b00,6'b000000,5'b00011,2'b01,5'b00001,6'b000011,3'b000};// ['ALU{A}->A', 'Flags']
MCODE0[1506]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1507]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1508]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1509]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1510]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1511]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// BD MOV SP, X
MCODE0[1512]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1513]={2'b10,2'b00,6'b000000,5'b00100,2'b00,5'b00000,6'b000000,3'b000};// ['X->SP']
MCODE0[1514]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1515]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1516]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1517]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1518]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1519]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// BE DAS
MCODE0[1520]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1521]={2'b00,2'b00,6'b000000,5'b00111,2'b01,5'b00000,6'b011111,3'b000};// ['ALU{A}->A', 'Flags']
MCODE0[1522]={2'b10,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[1523]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1524]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1525]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1526]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1527]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// BF MOV A, {X}+
MCODE0[1528]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1529]={2'b00,2'b00,6'b100101,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['X->AL', 'P->AH']
MCODE0[1530]={2'b00,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b000000,3'b000};// ['ALU{[AX]}->A', 'Flags']
MCODE0[1531]={2'b10,2'b00,6'b000000,5'b00000,2'b10,5'b00101,6'b000011,3'b000};// ['X++']
MCODE0[1532]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1533]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1534]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1535]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// C0 DI
MCODE0[1536]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1537]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[1538]={2'b10,2'b00,6'b000000,5'b01000,2'b00,5'b00000,6'b000000,3'b000};// ['Flags']
MCODE0[1539]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1540]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1541]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1542]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1543]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// C1 TCALL 12
MCODE0[1544]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1545]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[1546]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[1547]={2'b00,2'b10,6'b000000,5'b01101,2'b00,5'b00000,6'b000000,3'b101};// ['PCH->[SP]', 'SP--']
MCODE0[1548]={2'b00,2'b10,6'b000000,5'b01101,2'b00,5'b00000,6'b000000,3'b100};// ['PCL->[SP]', 'SP--']
MCODE0[1549]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[1550]={2'b00,2'b11,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['[VECT]->DR']
MCODE0[1551]={2'b10,2'b11,6'b000000,5'b01100,2'b00,5'b00000,6'b000000,3'b000};// ['[VECT]:DR->PC']
// C2 SET1 d.6
MCODE0[1552]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1553]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[1554]={2'b00,2'b01,6'b000000,5'b01011,2'b00,5'b10010,6'b010110,3'b000};// ['ALU{[AX]|40}', 'ALU{}->T']
MCODE0[1555]={2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001};// ['T->[AX]']
MCODE0[1556]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1557]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1558]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1559]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// C3 BBS d.6
MCODE0[1560]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1561]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[1562]={2'b00,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['[AX]->DR']
MCODE0[1563]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[1564]={2'b10,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->DR', 'PC++']
MCODE0[1565]={2'b00,2'b00,6'b000000,5'b01001,2'b00,5'b00000,6'b000000,3'b000};// ['PC+DR->PC']
MCODE0[1566]={2'b10,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[1567]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// C4 MOV d, A
MCODE0[1568]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1569]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[1570]={2'b00,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['[AX]']
MCODE0[1571]={2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b001};// ['A->[AX]']
MCODE0[1572]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1573]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1574]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1575]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// C5 MOV !a, A
MCODE0[1576]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1577]={2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'PC++']
MCODE0[1578]={2'b00,2'b00,6'b001000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AH', 'PC++']
MCODE0[1579]={2'b00,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['[AX]']
MCODE0[1580]={2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b001};// ['A->[AX]']
MCODE0[1581]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1582]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1583]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// C6 MOV {X}; A
MCODE0[1584]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1585]={2'b00,2'b00,6'b100101,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['X->AL', 'P->AH']
MCODE0[1586]={2'b00,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['[AX]']
MCODE0[1587]={2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b001};// ['A->[AX]']
MCODE0[1588]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1589]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1590]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1591]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// C7 MOV {d+X}; A
MCODE0[1592]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1593]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[1594]={2'b00,2'b00,6'b010000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['AL+X->AL']
MCODE0[1595]={2'b00,2'b01,6'b110000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['[AX]->DR', 'AL+1->AL']
MCODE0[1596]={2'b00,2'b01,6'b011010,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['[AX]->AH', 'DR->AL']
MCODE0[1597]={2'b00,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['[AX]']
MCODE0[1598]={2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b001};// ['A->[AX]']
MCODE0[1599]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// C8 CMP X, #i
MCODE0[1600]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1601]={2'b10,2'b00,6'b000000,5'b00010,2'b00,5'b00100,6'b010011,3'b000};// ['ALU{X-[PC]}', 'PC++', 'Flags']
MCODE0[1602]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1603]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1604]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1605]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1606]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1607]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// C9 MOV !a, X
MCODE0[1608]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1609]={2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'PC++']
MCODE0[1610]={2'b00,2'b00,6'b001000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AH', 'PC++']
MCODE0[1611]={2'b00,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['[AX]']
MCODE0[1612]={2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b00100,6'b000000,3'b001};// ['X->[AX]']
MCODE0[1613]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1614]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1615]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// CA MOV1 m.b, C
MCODE0[1616]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1617]={2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'PC++']
MCODE0[1618]={2'b00,2'b00,6'b001000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]&1F->AH', '[PC]->DR', 'PC++']
MCODE0[1619]={2'b00,2'b01,6'b000000,5'b01011,2'b00,5'b10010,6'b010101,3'b000};// ['ALU{[AX]}->T']
MCODE0[1620]={2'b00,2'b00,6'b000000,5'b01011,2'b00,5'b11111,6'b010110,3'b000};// ['ALU{T}->T']
MCODE0[1621]={2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001};// ['T->[AX]']
MCODE0[1622]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1623]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// CB MOV d, Y
MCODE0[1624]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1625]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[1626]={2'b00,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['[AX]']
MCODE0[1627]={2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01000,6'b000000,3'b001};// ['Y->[AX]']
MCODE0[1628]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1629]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1630]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1631]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// CC MOV !a, Y
MCODE0[1632]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1633]={2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'PC++']
MCODE0[1634]={2'b00,2'b00,6'b001000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AH', 'PC++']
MCODE0[1635]={2'b00,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['[AX]']
MCODE0[1636]={2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01000,6'b000000,3'b001};// ['Y->[AX]']
MCODE0[1637]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1638]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1639]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// CD MOV X, #i
MCODE0[1640]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1641]={2'b10,2'b00,6'b000000,5'b00010,2'b10,5'b00000,6'b000000,3'b000};// ['ALU{[PC]}->X', 'PC++', 'Flags']
MCODE0[1642]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1643]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1644]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1645]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1646]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1647]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// CE POP X
MCODE0[1648]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1649]={2'b00,2'b00,6'b000000,5'b10000,2'b00,5'b00000,6'b000000,3'b000};// ['SP++']
MCODE0[1650]={2'b00,2'b10,6'b000000,5'b00000,2'b10,5'b00000,6'b000000,3'b000};// ['[SP]->X']
MCODE0[1651]={2'b10,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[1652]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1653]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1654]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1655]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// CF MUL YA
MCODE0[1656]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1657]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b100000,3'b000};// ['ALU{Y*A}']
MCODE0[1658]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b100000,3'b000};// ['ALU{Y*A}']
MCODE0[1659]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b100000,3'b000};// ['ALU{Y*A}']
MCODE0[1660]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b100000,3'b000};// ['ALU{Y*A}']
MCODE0[1661]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b100000,3'b000};// ['ALU{Y*A}']
MCODE0[1662]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b100000,3'b000};// ['ALU{Y*A}']
MCODE0[1663]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b100000,3'b000};// ['ALU{Y*A}']
// D0 BNE
MCODE0[1664]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1665]={2'b10,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->DR', 'PC++']
MCODE0[1666]={2'b00,2'b00,6'b000000,5'b01001,2'b00,5'b00000,6'b000000,3'b000};// ['PC+DR->PC']
MCODE0[1667]={2'b10,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[1668]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1669]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1670]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1671]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// D1 TCALL 13
MCODE0[1672]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1673]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[1674]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[1675]={2'b00,2'b10,6'b000000,5'b01101,2'b00,5'b00000,6'b000000,3'b101};// ['PCH->[SP]', 'SP--']
MCODE0[1676]={2'b00,2'b10,6'b000000,5'b01101,2'b00,5'b00000,6'b000000,3'b100};// ['PCL->[SP]', 'SP--']
MCODE0[1677]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[1678]={2'b00,2'b11,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['[VECT]->DR']
MCODE0[1679]={2'b10,2'b11,6'b000000,5'b01100,2'b00,5'b00000,6'b000000,3'b000};// ['[VECT]:DR->PC']
// D2 CLR1 d.6
MCODE0[1680]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1681]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[1682]={2'b00,2'b01,6'b000000,5'b01011,2'b00,5'b10010,6'b010101,3'b000};// ['ALU{[AX]&~40}', 'ALU{}->T']
MCODE0[1683]={2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001};// ['T->[AX]']
MCODE0[1684]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1685]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1686]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1687]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// D3 BBC d.6
MCODE0[1688]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1689]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[1690]={2'b00,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['[AX]->DR']
MCODE0[1691]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[1692]={2'b10,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->DR', 'PC++']
MCODE0[1693]={2'b00,2'b00,6'b000000,5'b01001,2'b00,5'b00000,6'b000000,3'b000};// ['PC+DR->PC']
MCODE0[1694]={2'b10,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[1695]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// D4 MOV d+X, A
MCODE0[1696]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1697]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[1698]={2'b00,2'b00,6'b010000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['AL+X->AL']
MCODE0[1699]={2'b00,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['[AX]']
MCODE0[1700]={2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b001};// ['A->[AX]']
MCODE0[1701]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1702]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1703]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// D5 MOV !a+X, A
MCODE0[1704]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1705]={2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'PC++']
MCODE0[1706]={2'b00,2'b00,6'b011000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AH', 'AL+X->AL', 'PC++']
MCODE0[1707]={2'b00,2'b00,6'b001100,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['AH+Carry->AH']
MCODE0[1708]={2'b00,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['[AX]']
MCODE0[1709]={2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b001};// ['A->[AX]']
MCODE0[1710]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1711]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// D6 MOV !a+Y, A
MCODE0[1712]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1713]={2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'PC++']
MCODE0[1714]={2'b00,2'b00,6'b011001,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AH', 'AL+X->AL', 'PC++']
MCODE0[1715]={2'b00,2'b00,6'b001100,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['AH+Carry->AH']
MCODE0[1716]={2'b00,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['[AX]']
MCODE0[1717]={2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b001};// ['A->[AX]']
MCODE0[1718]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1719]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// D7 MOV {d}+Y, A
MCODE0[1720]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1721]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[1722]={2'b00,2'b01,6'b110000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['[AX]->DR', 'AL+1->AL']
MCODE0[1723]={2'b00,2'b01,6'b011011,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['[AX]->AH', 'DR+Y->AL']
MCODE0[1724]={2'b00,2'b00,6'b001100,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['AH+Carry->AH']
MCODE0[1725]={2'b00,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['[AX]']
MCODE0[1726]={2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b001};// ['A->[AX]']
MCODE0[1727]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// D8 MOV d, X
MCODE0[1728]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1729]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[1730]={2'b00,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['[AX]']
MCODE0[1731]={2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b00100,6'b000000,3'b001};// ['X->[AX]']
MCODE0[1732]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1733]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1734]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1735]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// D9 MOV d+Y, X
MCODE0[1736]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1737]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[1738]={2'b00,2'b00,6'b010001,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['AL+Y->AL']
MCODE0[1739]={2'b00,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['[AX]']
MCODE0[1740]={2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b00100,6'b000000,3'b001};// ['X->[AX]']
MCODE0[1741]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1742]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1743]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// DA MOV d, YA
MCODE0[1744]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1745]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[1746]={2'b00,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['[AX]']
MCODE0[1747]={2'b00,2'b01,6'b110000,5'b00000,2'b00,5'b00000,6'b000000,3'b001};// ['A->[AX]', 'AL+1->AL']
MCODE0[1748]={2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01000,6'b000000,3'b001};// ['Y->[AX]']
MCODE0[1749]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1750]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1751]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// DB MOV d+X, Y
MCODE0[1752]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1753]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[1754]={2'b00,2'b00,6'b010000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['AL+X->AL']
MCODE0[1755]={2'b00,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['[AX]']
MCODE0[1756]={2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01000,6'b000000,3'b001};// ['A->[AX]']
MCODE0[1757]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1758]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1759]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// DC DEC Y
MCODE0[1760]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1761]={2'b10,2'b00,6'b000000,5'b00011,2'b11,5'b01001,6'b000010,3'b000};// ['ALU{Y-1}', 'ALU{}->Y', 'Flags']
MCODE0[1762]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1763]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1764]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1765]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1766]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1767]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// DD MOV A, Y
MCODE0[1768]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1769]={2'b10,2'b00,6'b000000,5'b00011,2'b01,5'b01001,6'b000000,3'b000};// ['ALU{Y}->A', 'Flags']
MCODE0[1770]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1771]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1772]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1773]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1774]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1775]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// DE CBNE d+X, r
MCODE0[1776]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1777]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[1778]={2'b00,2'b00,6'b010000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['AL+X->AL']
MCODE0[1779]={2'b00,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b010011,3'b000};// ['ALU{[AX]}']
MCODE0[1780]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[1781]={2'b10,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->DR', 'PC++']
MCODE0[1782]={2'b00,2'b00,6'b000000,5'b01001,2'b00,5'b00000,6'b000000,3'b000};// ['PC+DR->PC']
MCODE0[1783]={2'b10,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
// DF DAA
MCODE0[1784]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1785]={2'b00,2'b00,6'b000000,5'b00111,2'b01,5'b00000,6'b011110,3'b000};// ['ALU{A}->A', 'Flags']
MCODE0[1786]={2'b10,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[1787]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1788]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1789]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1790]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1791]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// E0 CLRV
MCODE0[1792]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1793]={2'b10,2'b00,6'b000000,5'b01000,2'b00,5'b00000,6'b000000,3'b000};// ['Flags']
MCODE0[1794]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1795]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1796]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1797]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1798]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1799]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// E1 TCALL 14
MCODE0[1800]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1801]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[1802]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[1803]={2'b00,2'b10,6'b000000,5'b01101,2'b00,5'b00000,6'b000000,3'b101};// ['PCH->[SP]', 'SP--']
MCODE0[1804]={2'b00,2'b10,6'b000000,5'b01101,2'b00,5'b00000,6'b000000,3'b100};// ['PCL->[SP]', 'SP--']
MCODE0[1805]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[1806]={2'b00,2'b11,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['[VECT]->DR']
MCODE0[1807]={2'b10,2'b11,6'b000000,5'b01100,2'b00,5'b00000,6'b000000,3'b000};// ['[VECT]:DR->PC']
// E2 SET1 d.7
MCODE0[1808]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1809]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[1810]={2'b00,2'b01,6'b000000,5'b01011,2'b00,5'b10010,6'b010110,3'b000};// ['ALU{[AX]|80}', 'ALU{}->T']
MCODE0[1811]={2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001};// ['T->[AX]']
MCODE0[1812]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1813]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1814]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1815]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// E3 BBS d.7
MCODE0[1816]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1817]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[1818]={2'b00,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['[AX]->DR']
MCODE0[1819]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[1820]={2'b10,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->DR', 'PC++']
MCODE0[1821]={2'b00,2'b00,6'b000000,5'b01001,2'b00,5'b00000,6'b000000,3'b000};// ['PC+DR->PC']
MCODE0[1822]={2'b10,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[1823]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// E4 MOV A, d
MCODE0[1824]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1825]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[1826]={2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b000000,3'b000};// ['ALU{[AX]}->A', 'Flags']
MCODE0[1827]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1828]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1829]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1830]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1831]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// E5 MOV A, !a
MCODE0[1832]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1833]={2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'PC++']
MCODE0[1834]={2'b00,2'b00,6'b001000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AH', 'PC++']
MCODE0[1835]={2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b000000,3'b000};// ['ALU{[AX]}->A', 'Flags']
MCODE0[1836]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1837]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1838]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1839]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// E6 MOV A, {X}
MCODE0[1840]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1841]={2'b00,2'b00,6'b100101,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['X->AL', 'P->AH']
MCODE0[1842]={2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b000000,3'b000};// ['ALU{[AX]}->A', 'Flags']
MCODE0[1843]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1844]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1845]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1846]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1847]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// E7 MOV A, {d+X}
MCODE0[1848]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1849]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[1850]={2'b00,2'b00,6'b010000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['AL+X->AL']
MCODE0[1851]={2'b00,2'b01,6'b110000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['[AX]->DR', 'AL+1->AL']
MCODE0[1852]={2'b00,2'b01,6'b011010,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['[AX]->AH', 'DR->AL']
MCODE0[1853]={2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b000000,3'b000};// ['ALU{[AX]}->A', 'Flags']
MCODE0[1854]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1855]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// E8 MOV A, #i
MCODE0[1856]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1857]={2'b10,2'b00,6'b000000,5'b00010,2'b01,5'b00000,6'b000000,3'b000};// ['ALU{[PC]}->A', 'PC++', 'Flags']
MCODE0[1858]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1859]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1860]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1861]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1862]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1863]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// E9 X, !a
MCODE0[1864]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1865]={2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'PC++']
MCODE0[1866]={2'b00,2'b00,6'b001000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AH', 'PC++']
MCODE0[1867]={2'b10,2'b01,6'b000000,5'b00011,2'b10,5'b00000,6'b000000,3'b000};// ['ALU{[AX]}->X', 'Flags']
MCODE0[1868]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1869]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1870]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1871]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// EA NOT1 m.b
MCODE0[1872]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1873]={2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'PC++']
MCODE0[1874]={2'b00,2'b00,6'b001000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]&1F->AH', '[PC]->DR', 'PC++']
MCODE0[1875]={2'b00,2'b01,6'b000000,5'b01011,2'b00,5'b10010,6'b011011,3'b000};// ['ALU{[AX]}->T']
MCODE0[1876]={2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001};// ['T->[AX]']
MCODE0[1877]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1878]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1879]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// EB MOV Y, d
MCODE0[1880]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1881]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[1882]={2'b10,2'b01,6'b000000,5'b00011,2'b11,5'b00000,6'b000000,3'b000};// ['ALU{[AX]}->Y', 'Flags']
MCODE0[1883]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1884]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1885]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1886]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1887]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// EC Y, !a
MCODE0[1888]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1889]={2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'PC++']
MCODE0[1890]={2'b00,2'b00,6'b001000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AH', 'PC++']
MCODE0[1891]={2'b10,2'b01,6'b000000,5'b00011,2'b11,5'b00000,6'b000000,3'b000};// ['ALU{[AX]}->Y', 'Flags']
MCODE0[1892]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1893]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1894]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1895]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// ED NOT C
MCODE0[1896]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1897]={2'b00,2'b00,6'b000000,5'b01010,2'b00,5'b10100,6'b011100,3'b000};// ['C ^ 1']
MCODE0[1898]={2'b10,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[1899]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1900]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1901]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1902]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1903]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// EE POP Y
MCODE0[1904]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1905]={2'b00,2'b00,6'b000000,5'b10000,2'b00,5'b00000,6'b000000,3'b000};// ['SP++']
MCODE0[1906]={2'b00,2'b10,6'b000000,5'b00000,2'b11,5'b00000,6'b000000,3'b000};// ['[SP]->Y']
MCODE0[1907]={2'b10,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};//
MCODE0[1908]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1909]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1910]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1911]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// EF SLEEP
MCODE0[1912]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1913]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[1914]={2'b10,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[1915]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1916]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1917]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1918]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1919]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// F0 BEQ
MCODE0[1920]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1921]={2'b10,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->DR', 'PC++']
MCODE0[1922]={2'b00,2'b00,6'b000000,5'b01001,2'b00,5'b00000,6'b000000,3'b000};// ['PC+DR->PC']
MCODE0[1923]={2'b10,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[1924]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1925]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1926]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1927]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// F1 TCALL 15
MCODE0[1928]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1929]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[1930]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[1931]={2'b00,2'b10,6'b000000,5'b01101,2'b00,5'b00000,6'b000000,3'b101};// ['PCH->[SP]', 'SP--']
MCODE0[1932]={2'b00,2'b10,6'b000000,5'b01101,2'b00,5'b00000,6'b000000,3'b100};// ['PCL->[SP]', 'SP--']
MCODE0[1933]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[1934]={2'b00,2'b11,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['[VECT]->DR ']
MCODE0[1935]={2'b10,2'b11,6'b000000,5'b01100,2'b00,5'b00000,6'b000000,3'b000};// ['[VECT]:DR->PC ']
// F2 CLR1 d.7
MCODE0[1936]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1937]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[1938]={2'b00,2'b01,6'b000000,5'b01011,2'b00,5'b10010,6'b010101,3'b000};// ['ALU{[AX]&~80}', 'ALU{}->T']
MCODE0[1939]={2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001};// ['T->[AX]']
MCODE0[1940]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1941]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1942]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1943]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// F3 BBC d.7
MCODE0[1944]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1945]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[1946]={2'b00,2'b01,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['[AX]->DR']
MCODE0[1947]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[1948]={2'b10,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->DR', 'PC++']
MCODE0[1949]={2'b00,2'b00,6'b000000,5'b01001,2'b00,5'b00000,6'b000000,3'b000};// ['PC+DR->PC']
MCODE0[1950]={2'b10,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[1951]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// F4 MOV A, d+X
MCODE0[1952]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1953]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[1954]={2'b00,2'b00,6'b010000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['AL+X->AL']
MCODE0[1955]={2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b000000,3'b000};// ['ALU{[AX]}->A', 'Flags']
MCODE0[1956]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1957]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1958]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1959]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// F5 MOV A, !a+X
MCODE0[1960]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1961]={2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'PC++']
MCODE0[1962]={2'b00,2'b00,6'b011000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AH', 'AL+X->AL', 'PC++']
MCODE0[1963]={2'b00,2'b00,6'b001100,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['AH+Carry->AH']
MCODE0[1964]={2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b000000,3'b000};// ['ALU{[AX]}->A', 'Flags']
MCODE0[1965]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1966]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1967]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// F6 MOV A, !a+Y
MCODE0[1968]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1969]={2'b00,2'b00,6'b100000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'PC++']
MCODE0[1970]={2'b00,2'b00,6'b011001,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AH', 'AL+X->AL', 'PC++']
MCODE0[1971]={2'b00,2'b00,6'b001100,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['AH+Carry->AH']
MCODE0[1972]={2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b000000,3'b000};// ['ALU{[AX]}->A', 'Flags']
MCODE0[1973]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1974]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1975]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// F7 MOV A, {d}+Y
MCODE0[1976]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1977]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[1978]={2'b00,2'b01,6'b110000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['[AX]->DR', 'AL+1->AL']
MCODE0[1979]={2'b00,2'b01,6'b011011,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['[AX]->AH', 'DR+Y->AL']
MCODE0[1980]={2'b00,2'b00,6'b001100,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['AH+Carry->AH']
MCODE0[1981]={2'b10,2'b01,6'b000000,5'b00011,2'b01,5'b00000,6'b000000,3'b000};// ['ALU{[AX]}->A', 'Flags']
MCODE0[1982]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1983]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// F8 MOV X, d
MCODE0[1984]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1985]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[1986]={2'b10,2'b01,6'b000000,5'b00011,2'b10,5'b00000,6'b000000,3'b000};// ['ALU{[AX]}->X', 'Flags']
MCODE0[1987]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1988]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1989]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1990]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1991]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// F9 MOV X, d+Y
MCODE0[1992]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[1993]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[1994]={2'b00,2'b00,6'b010001,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['AL+Y->AL']
MCODE0[1995]={2'b10,2'b01,6'b000000,5'b00011,2'b10,5'b00000,6'b000000,3'b000};// ['ALU{[AX]}->X', 'Flags']
MCODE0[1996]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1997]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1998]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[1999]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// FA MOV dd, ds
MCODE0[2000]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[2001]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[2002]={2'b00,2'b01,6'b000000,5'b00110,2'b00,5'b00000,6'b000000,3'b000};// ['[AX]->T']
MCODE0[2003]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[2004]={2'b10,2'b01,6'b000000,5'b00000,2'b00,5'b01100,6'b000000,3'b001};// ['T->[AX]']
MCODE0[2005]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[2006]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[2007]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// FB MOV Y, d+X
MCODE0[2008]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[2009]={2'b00,2'b00,6'b100100,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->AL', 'P->AH', 'PC++']
MCODE0[2010]={2'b00,2'b00,6'b010000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// ['AL+X->AL']
MCODE0[2011]={2'b10,2'b01,6'b000000,5'b00011,2'b11,5'b00000,6'b000000,3'b000};// ['ALU{[AX]}->Y', 'Flags']
MCODE0[2012]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[2013]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[2014]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[2015]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// FC INC Y
MCODE0[2016]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[2017]={2'b10,2'b00,6'b000000,5'b00011,2'b11,5'b01001,6'b000011,3'b000};// ['ALU{Y}->Y', 'Flags']
MCODE0[2018]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[2019]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[2020]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[2021]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[2022]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[2023]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// FD MOV Y, A
MCODE0[2024]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[2025]={2'b10,2'b00,6'b000000,5'b00011,2'b11,5'b00001,6'b000000,3'b000};// ['ALU{A}->Y', 'Flags']
MCODE0[2026]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[2027]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[2028]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[2029]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[2030]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[2031]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// FE DBNZ Y, r
MCODE0[2032]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[2033]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[2034]={2'b00,2'b00,6'b000000,5'b00000,2'b11,5'b01001,6'b000010,3'b000};// ['ALU{Y}->Y', 'Flags']
MCODE0[2035]={2'b10,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['[PC]->DR', 'PC++']
MCODE0[2036]={2'b00,2'b00,6'b000000,5'b01001,2'b00,5'b00000,6'b000000,3'b000};// ['PC+DR->PC']
MCODE0[2037]={2'b10,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[2038]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[2039]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
// FF STOP
MCODE0[2040]={2'b00,2'b00,6'b000000,5'b00001,2'b00,5'b00000,6'b000000,3'b000};// ['PC++']
MCODE0[2041]={2'b00,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[2042]={2'b10,2'b00,6'b000000,5'b00000,2'b00,5'b00000,6'b000000,3'b000};// []
MCODE0[2043]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[2044]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[2045]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[2046]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
MCODE0[2047]={2'bXX,2'bXX,6'bXXXXXX,5'bXXXXX,2'bXX,5'bXXXXX,6'bXXXXXX,3'bXXX};
end
